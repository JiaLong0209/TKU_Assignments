
<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-32.95,39.6893,61.95,-63.2229</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>14.5,-13</position>
<gparam>LABEL_TEXT Go to https://cedar.to/vjyQw7 to download the latest version!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>14.5,-9.5</position>
<gparam>LABEL_TEXT Error: This file was made with a newer version of Cedar Logic!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 0>
</circuit>
<throw_away></throw_away>

	<version>2.3.8 | 2024-10-27 09:03:56</version><circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>444.834,-158.743,545.41,-212.241</PageViewport>
<gate>
<ID>368</ID>
<type>AA_LABEL</type>
<position>392,-151.5</position>
<gparam>LABEL_TEXT A4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>367</ID>
<type>AA_LABEL</type>
<position>392,-165</position>
<gparam>LABEL_TEXT A3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>366</ID>
<type>AA_LABEL</type>
<position>514,-274</position>
<gparam>LABEL_TEXT A5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>365</ID>
<type>AA_LABEL</type>
<position>514,-305</position>
<gparam>LABEL_TEXT B6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>164,-167</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>310</ID>
<type>AA_LABEL</type>
<position>514.5,-165</position>
<gparam>LABEL_TEXT A7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>164,-198</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>309</ID>
<type>DD_KEYPAD_HEX</type>
<position>522,-305</position>
<output>
<ID>OUT_0</ID>343 </output>
<output>
<ID>OUT_1</ID>349 </output>
<output>
<ID>OUT_2</ID>355 </output>
<output>
<ID>OUT_3</ID>361 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>51</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>296.5,-176</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>308</ID>
<type>AA_AND2</type>
<position>575.5,-274.5</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>352 </input>
<output>
<ID>OUT</ID>351 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>DD_KEYPAD_HEX</type>
<position>172,-166.5</position>
<output>
<ID>OUT_0</ID>25 </output>
<output>
<ID>OUT_1</ID>31 </output>
<output>
<ID>OUT_2</ID>37 </output>
<output>
<ID>OUT_3</ID>43 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>307</ID>
<type>AI_XOR2</type>
<position>561.5,-290.5</position>
<input>
<ID>IN_0</ID>347 </input>
<input>
<ID>IN_1</ID>346 </input>
<output>
<ID>OUT</ID>394 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>DD_KEYPAD_HEX</type>
<position>172,-211</position>
<output>
<ID>OUT_0</ID>26 </output>
<output>
<ID>OUT_1</ID>32 </output>
<output>
<ID>OUT_2</ID>38 </output>
<output>
<ID>OUT_3</ID>44 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>306</ID>
<type>AE_OR2</type>
<position>567.5,-280.5</position>
<input>
<ID>IN_0</ID>344 </input>
<input>
<ID>IN_1</ID>345 </input>
<output>
<ID>OUT</ID>352 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>AA_AND2</type>
<position>225.5,-219.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>305</ID>
<type>AI_XOR2</type>
<position>554,-284.5</position>
<input>
<ID>IN_0</ID>342 </input>
<input>
<ID>IN_1</ID>343 </input>
<output>
<ID>OUT</ID>347 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>47</ID>
<type>AI_XOR2</type>
<position>211.5,-235.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>304</ID>
<type>AA_AND2</type>
<position>561.5,-285.5</position>
<input>
<ID>IN_0</ID>347 </input>
<input>
<ID>IN_1</ID>346 </input>
<output>
<ID>OUT</ID>345 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AE_OR2</type>
<position>217.5,-225.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>AA_LABEL</type>
<position>514,-318</position>
<gparam>LABEL_TEXT B5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AI_XOR2</type>
<position>204,-229.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>302</ID>
<type>AE_OR2</type>
<position>581.5,-269.5</position>
<input>
<ID>IN_0</ID>350 </input>
<input>
<ID>IN_1</ID>351 </input>
<output>
<ID>OUT</ID>358 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AA_AND2</type>
<position>211.5,-230.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>301</ID>
<type>DD_KEYPAD_HEX</type>
<position>522,-260.5</position>
<output>
<ID>OUT_0</ID>342 </output>
<output>
<ID>OUT_1</ID>348 </output>
<output>
<ID>OUT_2</ID>354 </output>
<output>
<ID>OUT_3</ID>360 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>43</ID>
<type>AE_OR2</type>
<position>231.5,-214.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>300</ID>
<type>AA_AND2</type>
<position>554,-279.5</position>
<input>
<ID>IN_0</ID>342 </input>
<input>
<ID>IN_1</ID>343 </input>
<output>
<ID>OUT</ID>344 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>296.5,-185.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<input>
<ID>IN_2</ID>51 </input>
<input>
<ID>IN_3</ID>52 </input>
<input>
<ID>IN_4</ID>53 </input>
<input>
<ID>IN_5</ID>54 </input>
<input>
<ID>IN_6</ID>55 </input>
<input>
<ID>IN_7</ID>56 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>299</ID>
<type>AA_LABEL</type>
<position>514,-260.5</position>
<gparam>LABEL_TEXT A6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>DD_KEYPAD_HEX</type>
<position>172,-233.5</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>298</ID>
<type>AI_XOR2</type>
<position>568,-273.5</position>
<input>
<ID>IN_0</ID>348 </input>
<input>
<ID>IN_1</ID>349 </input>
<output>
<ID>OUT</ID>353 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>204,-224.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>297</ID>
<type>AI_XOR2</type>
<position>604.5,-254.5</position>
<input>
<ID>IN_0</ID>365 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>397 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>AI_XOR2</type>
<position>218,-218.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>296</ID>
<type>AI_XOR2</type>
<position>575.5,-279.5</position>
<input>
<ID>IN_0</ID>353 </input>
<input>
<ID>IN_1</ID>352 </input>
<output>
<ID>OUT</ID>395 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AI_XOR2</type>
<position>254.5,-199.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>295</ID>
<type>AA_AND2</type>
<position>597,-243.5</position>
<input>
<ID>IN_0</ID>360 </input>
<input>
<ID>IN_1</ID>361 </input>
<output>
<ID>OUT</ID>362 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AI_XOR2</type>
<position>225.5,-224.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>294</ID>
<type>AI_XOR2</type>
<position>597,-248.5</position>
<input>
<ID>IN_0</ID>360 </input>
<input>
<ID>IN_1</ID>361 </input>
<output>
<ID>OUT</ID>365 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>164.5,-233</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>293</ID>
<type>AA_AND2</type>
<position>582,-254.5</position>
<input>
<ID>IN_0</ID>354 </input>
<input>
<ID>IN_1</ID>355 </input>
<output>
<ID>OUT</ID>356 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_AND2</type>
<position>247,-188.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>292</ID>
<type>AA_AND2</type>
<position>589.5,-260.5</position>
<input>
<ID>IN_0</ID>359 </input>
<input>
<ID>IN_1</ID>358 </input>
<output>
<ID>OUT</ID>357 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>AI_XOR2</type>
<position>247,-193.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>291</ID>
<type>AE_OR2</type>
<position>595.5,-255.5</position>
<input>
<ID>IN_0</ID>356 </input>
<input>
<ID>IN_1</ID>357 </input>
<output>
<ID>OUT</ID>364 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AA_AND2</type>
<position>232,-199.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>290</ID>
<type>AA_AND2</type>
<position>568,-268.5</position>
<input>
<ID>IN_0</ID>348 </input>
<input>
<ID>IN_1</ID>349 </input>
<output>
<ID>OUT</ID>350 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_AND2</type>
<position>239.5,-205.5</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>289</ID>
<type>AE_OR2</type>
<position>610.5,-244.5</position>
<input>
<ID>IN_0</ID>362 </input>
<input>
<ID>IN_1</ID>363 </input>
<output>
<ID>OUT</ID>313 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AE_OR2</type>
<position>245.5,-200.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>288</ID>
<type>AA_AND2</type>
<position>604.5,-249.5</position>
<input>
<ID>IN_0</ID>365 </input>
<input>
<ID>IN_1</ID>364 </input>
<output>
<ID>OUT</ID>363 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_AND2</type>
<position>218,-213.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>287</ID>
<type>AI_XOR2</type>
<position>589.5,-265.5</position>
<input>
<ID>IN_0</ID>359 </input>
<input>
<ID>IN_1</ID>358 </input>
<output>
<ID>OUT</ID>396 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>AE_OR2</type>
<position>260.5,-189.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>286</ID>
<type>AI_XOR2</type>
<position>582,-259.5</position>
<input>
<ID>IN_0</ID>354 </input>
<input>
<ID>IN_1</ID>355 </input>
<output>
<ID>OUT</ID>359 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_AND2</type>
<position>254.5,-194.5</position>
<input>
<ID>IN_0</ID>48 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>285</ID>
<type>AI_XOR2</type>
<position>582,-311.5</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>383 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>AI_XOR2</type>
<position>239.5,-210.5</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>284</ID>
<type>AI_XOR2</type>
<position>589.5,-317.5</position>
<input>
<ID>IN_0</ID>383 </input>
<input>
<ID>IN_1</ID>382 </input>
<output>
<ID>OUT</ID>392 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AI_XOR2</type>
<position>232,-204.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>283</ID>
<type>AA_AND2</type>
<position>604.5,-301.5</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>388 </input>
<output>
<ID>OUT</ID>387 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AI_XOR2</type>
<position>232,-152.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>282</ID>
<type>AE_OR2</type>
<position>610.5,-296.5</position>
<input>
<ID>IN_0</ID>386 </input>
<input>
<ID>IN_1</ID>387 </input>
<output>
<ID>OUT</ID>346 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AI_XOR2</type>
<position>239.5,-158.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>281</ID>
<type>AA_AND2</type>
<position>568,-320.5</position>
<input>
<ID>IN_0</ID>372 </input>
<input>
<ID>IN_1</ID>373 </input>
<output>
<ID>OUT</ID>374 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_AND2</type>
<position>254.5,-142.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>280</ID>
<type>AE_OR2</type>
<position>595.5,-307.5</position>
<input>
<ID>IN_0</ID>380 </input>
<input>
<ID>IN_1</ID>381 </input>
<output>
<ID>OUT</ID>388 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AE_OR2</type>
<position>260.5,-137.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>279</ID>
<type>AA_AND2</type>
<position>589.5,-312.5</position>
<input>
<ID>IN_0</ID>383 </input>
<input>
<ID>IN_1</ID>382 </input>
<output>
<ID>OUT</ID>381 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_AND2</type>
<position>218,-161.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>278</ID>
<type>AA_AND2</type>
<position>582,-306.5</position>
<input>
<ID>IN_0</ID>378 </input>
<input>
<ID>IN_1</ID>379 </input>
<output>
<ID>OUT</ID>380 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_OR2</type>
<position>245.5,-148.5</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>277</ID>
<type>AI_XOR2</type>
<position>597,-300.5</position>
<input>
<ID>IN_0</ID>384 </input>
<input>
<ID>IN_1</ID>385 </input>
<output>
<ID>OUT</ID>389 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AA_AND2</type>
<position>239.5,-153.5</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>276</ID>
<type>AA_AND2</type>
<position>597,-295.5</position>
<input>
<ID>IN_0</ID>384 </input>
<input>
<ID>IN_1</ID>385 </input>
<output>
<ID>OUT</ID>386 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>232,-147.5</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AI_XOR2</type>
<position>247,-141.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>274</ID>
<type>AI_XOR2</type>
<position>575.5,-331.5</position>
<input>
<ID>IN_0</ID>377 </input>
<input>
<ID>IN_1</ID>376 </input>
<output>
<ID>OUT</ID>391 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AA_AND2</type>
<position>247,-136.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>273</ID>
<type>AI_XOR2</type>
<position>604.5,-306.5</position>
<input>
<ID>IN_0</ID>389 </input>
<input>
<ID>IN_1</ID>388 </input>
<output>
<ID>OUT</ID>393 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AI_XOR2</type>
<position>225.5,-172.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>54 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>272</ID>
<type>AI_XOR2</type>
<position>568,-325.5</position>
<input>
<ID>IN_0</ID>372 </input>
<input>
<ID>IN_1</ID>373 </input>
<output>
<ID>OUT</ID>377 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AI_XOR2</type>
<position>254.5,-147.5</position>
<input>
<ID>IN_0</ID>24 </input>
<input>
<ID>IN_1</ID>23 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>271</ID>
<type>AA_AND2</type>
<position>554,-331.5</position>
<input>
<ID>IN_0</ID>366 </input>
<input>
<ID>IN_1</ID>367 </input>
<output>
<ID>OUT</ID>368 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>AI_XOR2</type>
<position>218,-166.5</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>164,-153.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>269</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>646.5,-292.5</position>
<input>
<ID>IN_0</ID>390 </input>
<input>
<ID>IN_1</ID>391 </input>
<input>
<ID>IN_2</ID>392 </input>
<input>
<ID>IN_3</ID>393 </input>
<input>
<ID>IN_4</ID>394 </input>
<input>
<ID>IN_5</ID>395 </input>
<input>
<ID>IN_6</ID>396 </input>
<input>
<ID>IN_7</ID>397 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_AND2</type>
<position>204,-172.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>268</ID>
<type>AE_OR2</type>
<position>581.5,-321.5</position>
<input>
<ID>IN_0</ID>374 </input>
<input>
<ID>IN_1</ID>375 </input>
<output>
<ID>OUT</ID>382 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>222.5,-131.5</position>
<gparam>LABEL_TEXT 8-Bits Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>267</ID>
<type>AA_AND2</type>
<position>561.5,-337.5</position>
<input>
<ID>IN_0</ID>371 </input>
<input>
<ID>IN_1</ID>370 </input>
<output>
<ID>OUT</ID>369 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>DD_KEYPAD_HEX</type>
<position>172,-153.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<output>
<ID>OUT_1</ID>7 </output>
<output>
<ID>OUT_2</ID>13 </output>
<output>
<ID>OUT_3</ID>19 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>266</ID>
<type>AI_XOR2</type>
<position>554,-336.5</position>
<input>
<ID>IN_0</ID>366 </input>
<input>
<ID>IN_1</ID>367 </input>
<output>
<ID>OUT</ID>371 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AE_OR2</type>
<position>231.5,-162.5</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>265</ID>
<type>AE_OR2</type>
<position>567.5,-332.5</position>
<input>
<ID>IN_0</ID>368 </input>
<input>
<ID>IN_1</ID>369 </input>
<output>
<ID>OUT</ID>376 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>164,-211</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>264</ID>
<type>AI_XOR2</type>
<position>561.5,-342.5</position>
<input>
<ID>IN_0</ID>371 </input>
<input>
<ID>IN_1</ID>370 </input>
<output>
<ID>OUT</ID>390 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND2</type>
<position>211.5,-178.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>263</ID>
<type>AA_LABEL</type>
<position>391,-274</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AI_XOR2</type>
<position>204,-177.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>262</ID>
<type>AA_LABEL</type>
<position>391,-305</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AE_OR2</type>
<position>217.5,-173.5</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>3</ID>
<type>AI_XOR2</type>
<position>211.5,-183.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>260</ID>
<type>DD_KEYPAD_HEX</type>
<position>399,-273.5</position>
<output>
<ID>OUT_0</ID>252 </output>
<output>
<ID>OUT_1</ID>258 </output>
<output>
<ID>OUT_2</ID>264 </output>
<output>
<ID>OUT_3</ID>270 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>2</ID>
<type>AA_AND2</type>
<position>225.5,-167.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>10 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>259</ID>
<type>DD_KEYPAD_HEX</type>
<position>399,-318</position>
<output>
<ID>OUT_0</ID>253 </output>
<output>
<ID>OUT_1</ID>259 </output>
<output>
<ID>OUT_2</ID>265 </output>
<output>
<ID>OUT_3</ID>271 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>1</ID>
<type>DD_KEYPAD_HEX</type>
<position>172,-198</position>
<output>
<ID>OUT_0</ID>2 </output>
<output>
<ID>OUT_1</ID>8 </output>
<output>
<ID>OUT_2</ID>14 </output>
<output>
<ID>OUT_3</ID>20 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_AND2</type>
<position>452.5,-326.5</position>
<input>
<ID>IN_0</ID>263 </input>
<input>
<ID>IN_1</ID>262 </input>
<output>
<ID>OUT</ID>261 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>158</ID>
<type>DD_KEYPAD_HEX</type>
<position>399.5,-196</position>
<output>
<ID>OUT_0</ID>172 </output>
<output>
<ID>OUT_1</ID>178 </output>
<output>
<ID>OUT_2</ID>184 </output>
<output>
<ID>OUT_3</ID>190 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_AND2</type>
<position>453,-165.5</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>180 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>AI_XOR2</type>
<position>439,-181.5</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>175 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>AE_OR2</type>
<position>445,-171.5</position>
<input>
<ID>IN_0</ID>173 </input>
<input>
<ID>IN_1</ID>174 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>AI_XOR2</type>
<position>431.5,-175.5</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>163</ID>
<type>AA_AND2</type>
<position>439,-176.5</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>175 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_LABEL</type>
<position>391.5,-209</position>
<gparam>LABEL_TEXT B3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>165</ID>
<type>AE_OR2</type>
<position>459,-160.5</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>180 </input>
<output>
<ID>OUT</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>DD_KEYPAD_HEX</type>
<position>399.5,-151.5</position>
<output>
<ID>OUT_0</ID>171 </output>
<output>
<ID>OUT_1</ID>177 </output>
<output>
<ID>OUT_2</ID>183 </output>
<output>
<ID>OUT_3</ID>189 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>167</ID>
<type>AA_LABEL</type>
<position>450,-129.5</position>
<gparam>LABEL_TEXT 8-Bits Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_AND2</type>
<position>431.5,-170.5</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AI_XOR2</type>
<position>445.5,-164.5</position>
<input>
<ID>IN_0</ID>177 </input>
<input>
<ID>IN_1</ID>178 </input>
<output>
<ID>OUT</ID>182 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>AI_XOR2</type>
<position>482,-145.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>193 </input>
<output>
<ID>OUT</ID>226 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>AI_XOR2</type>
<position>453,-170.5</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_AND2</type>
<position>474.5,-134.5</position>
<input>
<ID>IN_0</ID>189 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>191 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>174</ID>
<type>AI_XOR2</type>
<position>474.5,-139.5</position>
<input>
<ID>IN_0</ID>189 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_AND2</type>
<position>459.5,-145.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>184 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>176</ID>
<type>AA_AND2</type>
<position>467,-151.5</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>186 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>AE_OR2</type>
<position>473,-146.5</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>186 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>178</ID>
<type>AA_AND2</type>
<position>445.5,-159.5</position>
<input>
<ID>IN_0</ID>177 </input>
<input>
<ID>IN_1</ID>178 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>AE_OR2</type>
<position>488,-135.5</position>
<input>
<ID>IN_0</ID>191 </input>
<input>
<ID>IN_1</ID>192 </input>
<output>
<ID>OUT</ID>370 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>AA_AND2</type>
<position>482,-140.5</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>193 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>181</ID>
<type>AI_XOR2</type>
<position>467,-156.5</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>182</ID>
<type>AI_XOR2</type>
<position>459.5,-150.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>184 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>AI_XOR2</type>
<position>459.5,-202.5</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>212 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>184</ID>
<type>AI_XOR2</type>
<position>467,-208.5</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>185</ID>
<type>AA_AND2</type>
<position>482,-192.5</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>186</ID>
<type>AE_OR2</type>
<position>488,-187.5</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>216 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_AND2</type>
<position>445.5,-211.5</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>202 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>AE_OR2</type>
<position>473,-198.5</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>210 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>189</ID>
<type>AA_AND2</type>
<position>467,-203.5</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>190</ID>
<type>AA_AND2</type>
<position>459.5,-197.5</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>191</ID>
<type>AI_XOR2</type>
<position>474.5,-191.5</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>218 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_AND2</type>
<position>474.5,-186.5</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>194</ID>
<type>AI_XOR2</type>
<position>453,-222.5</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>205 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>195</ID>
<type>AI_XOR2</type>
<position>482,-197.5</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>AI_XOR2</type>
<position>445.5,-216.5</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>202 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_AND2</type>
<position>431.5,-222.5</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>196 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>505.5,-184</position>
<input>
<ID>IN_0</ID>219 </input>
<input>
<ID>IN_1</ID>220 </input>
<input>
<ID>IN_2</ID>221 </input>
<input>
<ID>IN_3</ID>222 </input>
<input>
<ID>IN_4</ID>223 </input>
<input>
<ID>IN_6</ID>225 </input>
<input>
<ID>IN_7</ID>226 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 223</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>200</ID>
<type>AE_OR2</type>
<position>459,-212.5</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>204 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>AA_AND2</type>
<position>439,-228.5</position>
<input>
<ID>IN_0</ID>200 </input>
<input>
<ID>IN_1</ID>199 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>AI_XOR2</type>
<position>431.5,-227.5</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>196 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>203</ID>
<type>AE_OR2</type>
<position>445,-223.5</position>
<input>
<ID>IN_0</ID>197 </input>
<input>
<ID>IN_1</ID>198 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>204</ID>
<type>AI_XOR2</type>
<position>439,-233.5</position>
<input>
<ID>IN_0</ID>200 </input>
<input>
<ID>IN_1</ID>199 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>AA_AND2</type>
<position>453,-217.5</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>205 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>206</ID>
<type>DD_KEYPAD_HEX</type>
<position>399.5,-209</position>
<output>
<ID>OUT_0</ID>196 </output>
<output>
<ID>OUT_1</ID>202 </output>
<output>
<ID>OUT_2</ID>208 </output>
<output>
<ID>OUT_3</ID>214 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>207</ID>
<type>DD_KEYPAD_HEX</type>
<position>399.5,-164.5</position>
<output>
<ID>OUT_0</ID>195 </output>
<output>
<ID>OUT_1</ID>201 </output>
<output>
<ID>OUT_2</ID>207 </output>
<output>
<ID>OUT_3</ID>213 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_LABEL</type>
<position>391.5,-196</position>
<gparam>LABEL_TEXT B4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>DD_KEYPAD_HEX</type>
<position>399,-305</position>
<output>
<ID>OUT_0</ID>229 </output>
<output>
<ID>OUT_1</ID>235 </output>
<output>
<ID>OUT_2</ID>241 </output>
<output>
<ID>OUT_3</ID>247 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_AND2</type>
<position>452.5,-274.5</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>237 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>AI_XOR2</type>
<position>438.5,-290.5</position>
<input>
<ID>IN_0</ID>233 </input>
<input>
<ID>IN_1</ID>232 </input>
<output>
<ID>OUT</ID>280 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>214</ID>
<type>AE_OR2</type>
<position>444.5,-280.5</position>
<input>
<ID>IN_0</ID>230 </input>
<input>
<ID>IN_1</ID>231 </input>
<output>
<ID>OUT</ID>238 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AI_XOR2</type>
<position>431,-284.5</position>
<input>
<ID>IN_0</ID>228 </input>
<input>
<ID>IN_1</ID>229 </input>
<output>
<ID>OUT</ID>233 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_AND2</type>
<position>438.5,-285.5</position>
<input>
<ID>IN_0</ID>233 </input>
<input>
<ID>IN_1</ID>232 </input>
<output>
<ID>OUT</ID>231 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>391,-318</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>AE_OR2</type>
<position>458.5,-269.5</position>
<input>
<ID>IN_0</ID>236 </input>
<input>
<ID>IN_1</ID>237 </input>
<output>
<ID>OUT</ID>244 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>219</ID>
<type>DD_KEYPAD_HEX</type>
<position>399,-260.5</position>
<output>
<ID>OUT_0</ID>228 </output>
<output>
<ID>OUT_1</ID>234 </output>
<output>
<ID>OUT_2</ID>240 </output>
<output>
<ID>OUT_3</ID>246 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>431,-279.5</position>
<input>
<ID>IN_0</ID>228 </input>
<input>
<ID>IN_1</ID>229 </input>
<output>
<ID>OUT</ID>230 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>391,-260.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>223</ID>
<type>AI_XOR2</type>
<position>445,-273.5</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>235 </input>
<output>
<ID>OUT</ID>239 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>224</ID>
<type>AI_XOR2</type>
<position>481.5,-254.5</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>250 </input>
<output>
<ID>OUT</ID>283 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>AI_XOR2</type>
<position>452.5,-279.5</position>
<input>
<ID>IN_0</ID>239 </input>
<input>
<ID>IN_1</ID>238 </input>
<output>
<ID>OUT</ID>281 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>226</ID>
<type>AA_AND2</type>
<position>474,-243.5</position>
<input>
<ID>IN_0</ID>246 </input>
<input>
<ID>IN_1</ID>247 </input>
<output>
<ID>OUT</ID>248 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>AI_XOR2</type>
<position>474,-248.5</position>
<input>
<ID>IN_0</ID>246 </input>
<input>
<ID>IN_1</ID>247 </input>
<output>
<ID>OUT</ID>251 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AA_AND2</type>
<position>459,-254.5</position>
<input>
<ID>IN_0</ID>240 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>242 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>229</ID>
<type>AA_AND2</type>
<position>466.5,-260.5</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>243 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>AE_OR2</type>
<position>472.5,-255.5</position>
<input>
<ID>IN_0</ID>242 </input>
<input>
<ID>IN_1</ID>243 </input>
<output>
<ID>OUT</ID>250 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>231</ID>
<type>AA_AND2</type>
<position>445,-268.5</position>
<input>
<ID>IN_0</ID>234 </input>
<input>
<ID>IN_1</ID>235 </input>
<output>
<ID>OUT</ID>236 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>232</ID>
<type>AE_OR2</type>
<position>487.5,-244.5</position>
<input>
<ID>IN_0</ID>248 </input>
<input>
<ID>IN_1</ID>249 </input>
<output>
<ID>OUT</ID>199 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_AND2</type>
<position>481.5,-249.5</position>
<input>
<ID>IN_0</ID>251 </input>
<input>
<ID>IN_1</ID>250 </input>
<output>
<ID>OUT</ID>249 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>234</ID>
<type>AI_XOR2</type>
<position>466.5,-265.5</position>
<input>
<ID>IN_0</ID>245 </input>
<input>
<ID>IN_1</ID>244 </input>
<output>
<ID>OUT</ID>282 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>235</ID>
<type>AI_XOR2</type>
<position>459,-259.5</position>
<input>
<ID>IN_0</ID>240 </input>
<input>
<ID>IN_1</ID>241 </input>
<output>
<ID>OUT</ID>245 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>236</ID>
<type>AI_XOR2</type>
<position>459,-311.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>269 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>237</ID>
<type>AI_XOR2</type>
<position>466.5,-317.5</position>
<input>
<ID>IN_0</ID>269 </input>
<input>
<ID>IN_1</ID>268 </input>
<output>
<ID>OUT</ID>278 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>238</ID>
<type>AA_AND2</type>
<position>481.5,-301.5</position>
<input>
<ID>IN_0</ID>275 </input>
<input>
<ID>IN_1</ID>274 </input>
<output>
<ID>OUT</ID>273 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>239</ID>
<type>AE_OR2</type>
<position>487.5,-296.5</position>
<input>
<ID>IN_0</ID>272 </input>
<input>
<ID>IN_1</ID>273 </input>
<output>
<ID>OUT</ID>232 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>AA_AND2</type>
<position>445,-320.5</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>259 </input>
<output>
<ID>OUT</ID>260 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>241</ID>
<type>AE_OR2</type>
<position>472.5,-307.5</position>
<input>
<ID>IN_0</ID>266 </input>
<input>
<ID>IN_1</ID>267 </input>
<output>
<ID>OUT</ID>274 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>242</ID>
<type>AA_AND2</type>
<position>466.5,-312.5</position>
<input>
<ID>IN_0</ID>269 </input>
<input>
<ID>IN_1</ID>268 </input>
<output>
<ID>OUT</ID>267 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>243</ID>
<type>AA_AND2</type>
<position>459,-306.5</position>
<input>
<ID>IN_0</ID>264 </input>
<input>
<ID>IN_1</ID>265 </input>
<output>
<ID>OUT</ID>266 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>244</ID>
<type>AI_XOR2</type>
<position>474,-300.5</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>271 </input>
<output>
<ID>OUT</ID>275 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>245</ID>
<type>AA_AND2</type>
<position>474,-295.5</position>
<input>
<ID>IN_0</ID>270 </input>
<input>
<ID>IN_1</ID>271 </input>
<output>
<ID>OUT</ID>272 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>246</ID>
<type>AA_LABEL</type>
<position>391.5,-340</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>247</ID>
<type>AI_XOR2</type>
<position>452.5,-331.5</position>
<input>
<ID>IN_0</ID>263 </input>
<input>
<ID>IN_1</ID>262 </input>
<output>
<ID>OUT</ID>277 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>AI_XOR2</type>
<position>481.5,-306.5</position>
<input>
<ID>IN_0</ID>275 </input>
<input>
<ID>IN_1</ID>274 </input>
<output>
<ID>OUT</ID>279 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>249</ID>
<type>AI_XOR2</type>
<position>445,-325.5</position>
<input>
<ID>IN_0</ID>258 </input>
<input>
<ID>IN_1</ID>259 </input>
<output>
<ID>OUT</ID>263 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>250</ID>
<type>AA_AND2</type>
<position>431,-331.5</position>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>253 </input>
<output>
<ID>OUT</ID>254 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>251</ID>
<type>DD_KEYPAD_HEX</type>
<position>399,-340.5</position>
<output>
<ID>OUT_0</ID>256 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>252</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>503.5,-292.5</position>
<input>
<ID>IN_0</ID>276 </input>
<input>
<ID>IN_1</ID>277 </input>
<input>
<ID>IN_2</ID>278 </input>
<input>
<ID>IN_3</ID>279 </input>
<input>
<ID>IN_4</ID>280 </input>
<input>
<ID>IN_5</ID>281 </input>
<input>
<ID>IN_6</ID>282 </input>
<input>
<ID>IN_7</ID>283 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>253</ID>
<type>AE_OR2</type>
<position>458.5,-321.5</position>
<input>
<ID>IN_0</ID>260 </input>
<input>
<ID>IN_1</ID>261 </input>
<output>
<ID>OUT</ID>268 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_AND2</type>
<position>438.5,-337.5</position>
<input>
<ID>IN_0</ID>257 </input>
<input>
<ID>IN_1</ID>256 </input>
<output>
<ID>OUT</ID>255 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>255</ID>
<type>AI_XOR2</type>
<position>431,-336.5</position>
<input>
<ID>IN_0</ID>252 </input>
<input>
<ID>IN_1</ID>253 </input>
<output>
<ID>OUT</ID>257 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>256</ID>
<type>AE_OR2</type>
<position>444.5,-332.5</position>
<input>
<ID>IN_0</ID>254 </input>
<input>
<ID>IN_1</ID>255 </input>
<output>
<ID>OUT</ID>262 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>257</ID>
<type>AI_XOR2</type>
<position>438.5,-342.5</position>
<input>
<ID>IN_0</ID>257 </input>
<input>
<ID>IN_1</ID>256 </input>
<output>
<ID>OUT</ID>276 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>311</ID>
<type>AA_LABEL</type>
<position>514.5,-196</position>
<gparam>LABEL_TEXT B8</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>312</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>647,-174</position>
<input>
<ID>IN_0</ID>341 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>313</ID>
<type>DD_KEYPAD_HEX</type>
<position>522.5,-164.5</position>
<output>
<ID>OUT_0</ID>309 </output>
<output>
<ID>OUT_1</ID>315 </output>
<output>
<ID>OUT_2</ID>321 </output>
<output>
<ID>OUT_3</ID>327 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>314</ID>
<type>DD_KEYPAD_HEX</type>
<position>522.5,-209</position>
<output>
<ID>OUT_0</ID>310 </output>
<output>
<ID>OUT_1</ID>316 </output>
<output>
<ID>OUT_2</ID>322 </output>
<output>
<ID>OUT_3</ID>328 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>315</ID>
<type>AA_AND2</type>
<position>576,-217.5</position>
<input>
<ID>IN_0</ID>320 </input>
<input>
<ID>IN_1</ID>319 </input>
<output>
<ID>OUT</ID>318 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>316</ID>
<type>AI_XOR2</type>
<position>562,-233.5</position>
<input>
<ID>IN_0</ID>314 </input>
<input>
<ID>IN_1</ID>313 </input>
<output>
<ID>OUT</ID>333 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>317</ID>
<type>AE_OR2</type>
<position>568,-223.5</position>
<input>
<ID>IN_0</ID>311 </input>
<input>
<ID>IN_1</ID>312 </input>
<output>
<ID>OUT</ID>319 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>318</ID>
<type>AI_XOR2</type>
<position>554.5,-227.5</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>310 </input>
<output>
<ID>OUT</ID>314 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>319</ID>
<type>AA_AND2</type>
<position>562,-228.5</position>
<input>
<ID>IN_0</ID>314 </input>
<input>
<ID>IN_1</ID>313 </input>
<output>
<ID>OUT</ID>312 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>320</ID>
<type>AE_OR2</type>
<position>582,-212.5</position>
<input>
<ID>IN_0</ID>317 </input>
<input>
<ID>IN_1</ID>318 </input>
<output>
<ID>OUT</ID>325 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>321</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>647,-183.5</position>
<input>
<ID>IN_0</ID>333 </input>
<input>
<ID>IN_1</ID>334 </input>
<input>
<ID>IN_2</ID>335 </input>
<input>
<ID>IN_3</ID>336 </input>
<input>
<ID>IN_4</ID>337 </input>
<input>
<ID>IN_5</ID>338 </input>
<input>
<ID>IN_6</ID>339 </input>
<input>
<ID>IN_7</ID>340 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>322</ID>
<type>AA_AND2</type>
<position>554.5,-222.5</position>
<input>
<ID>IN_0</ID>309 </input>
<input>
<ID>IN_1</ID>310 </input>
<output>
<ID>OUT</ID>311 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>323</ID>
<type>AI_XOR2</type>
<position>568.5,-216.5</position>
<input>
<ID>IN_0</ID>315 </input>
<input>
<ID>IN_1</ID>316 </input>
<output>
<ID>OUT</ID>320 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>324</ID>
<type>AI_XOR2</type>
<position>605,-197.5</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>331 </input>
<output>
<ID>OUT</ID>336 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>325</ID>
<type>AI_XOR2</type>
<position>576,-222.5</position>
<input>
<ID>IN_0</ID>320 </input>
<input>
<ID>IN_1</ID>319 </input>
<output>
<ID>OUT</ID>334 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>326</ID>
<type>AA_AND2</type>
<position>597.5,-186.5</position>
<input>
<ID>IN_0</ID>327 </input>
<input>
<ID>IN_1</ID>328 </input>
<output>
<ID>OUT</ID>329 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>327</ID>
<type>AI_XOR2</type>
<position>597.5,-191.5</position>
<input>
<ID>IN_0</ID>327 </input>
<input>
<ID>IN_1</ID>328 </input>
<output>
<ID>OUT</ID>332 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>328</ID>
<type>AA_AND2</type>
<position>582.5,-197.5</position>
<input>
<ID>IN_0</ID>321 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>323 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>329</ID>
<type>AA_AND2</type>
<position>590,-203.5</position>
<input>
<ID>IN_0</ID>326 </input>
<input>
<ID>IN_1</ID>325 </input>
<output>
<ID>OUT</ID>324 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>330</ID>
<type>AE_OR2</type>
<position>596,-198.5</position>
<input>
<ID>IN_0</ID>323 </input>
<input>
<ID>IN_1</ID>324 </input>
<output>
<ID>OUT</ID>331 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>331</ID>
<type>AA_AND2</type>
<position>568.5,-211.5</position>
<input>
<ID>IN_0</ID>315 </input>
<input>
<ID>IN_1</ID>316 </input>
<output>
<ID>OUT</ID>317 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>332</ID>
<type>AE_OR2</type>
<position>611,-187.5</position>
<input>
<ID>IN_0</ID>329 </input>
<input>
<ID>IN_1</ID>330 </input>
<output>
<ID>OUT</ID>289 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>333</ID>
<type>AA_AND2</type>
<position>605,-192.5</position>
<input>
<ID>IN_0</ID>332 </input>
<input>
<ID>IN_1</ID>331 </input>
<output>
<ID>OUT</ID>330 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>334</ID>
<type>AI_XOR2</type>
<position>590,-208.5</position>
<input>
<ID>IN_0</ID>326 </input>
<input>
<ID>IN_1</ID>325 </input>
<output>
<ID>OUT</ID>335 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>335</ID>
<type>AI_XOR2</type>
<position>582.5,-202.5</position>
<input>
<ID>IN_0</ID>321 </input>
<input>
<ID>IN_1</ID>322 </input>
<output>
<ID>OUT</ID>326 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>336</ID>
<type>AI_XOR2</type>
<position>582.5,-150.5</position>
<input>
<ID>IN_0</ID>297 </input>
<input>
<ID>IN_1</ID>298 </input>
<output>
<ID>OUT</ID>302 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>337</ID>
<type>AI_XOR2</type>
<position>590,-156.5</position>
<input>
<ID>IN_0</ID>302 </input>
<input>
<ID>IN_1</ID>301 </input>
<output>
<ID>OUT</ID>339 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>338</ID>
<type>AA_AND2</type>
<position>605,-140.5</position>
<input>
<ID>IN_0</ID>308 </input>
<input>
<ID>IN_1</ID>307 </input>
<output>
<ID>OUT</ID>306 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>339</ID>
<type>AE_OR2</type>
<position>611,-135.5</position>
<input>
<ID>IN_0</ID>305 </input>
<input>
<ID>IN_1</ID>306 </input>
<output>
<ID>OUT</ID>341 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>340</ID>
<type>AA_AND2</type>
<position>568.5,-159.5</position>
<input>
<ID>IN_0</ID>291 </input>
<input>
<ID>IN_1</ID>292 </input>
<output>
<ID>OUT</ID>293 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>341</ID>
<type>AE_OR2</type>
<position>596,-146.5</position>
<input>
<ID>IN_0</ID>299 </input>
<input>
<ID>IN_1</ID>300 </input>
<output>
<ID>OUT</ID>307 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>342</ID>
<type>AA_AND2</type>
<position>590,-151.5</position>
<input>
<ID>IN_0</ID>302 </input>
<input>
<ID>IN_1</ID>301 </input>
<output>
<ID>OUT</ID>300 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>343</ID>
<type>AA_AND2</type>
<position>582.5,-145.5</position>
<input>
<ID>IN_0</ID>297 </input>
<input>
<ID>IN_1</ID>298 </input>
<output>
<ID>OUT</ID>299 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>344</ID>
<type>AI_XOR2</type>
<position>597.5,-139.5</position>
<input>
<ID>IN_0</ID>303 </input>
<input>
<ID>IN_1</ID>304 </input>
<output>
<ID>OUT</ID>308 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>345</ID>
<type>AA_AND2</type>
<position>597.5,-134.5</position>
<input>
<ID>IN_0</ID>303 </input>
<input>
<ID>IN_1</ID>304 </input>
<output>
<ID>OUT</ID>305 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>346</ID>
<type>AI_XOR2</type>
<position>576,-170.5</position>
<input>
<ID>IN_0</ID>296 </input>
<input>
<ID>IN_1</ID>295 </input>
<output>
<ID>OUT</ID>338 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>347</ID>
<type>AI_XOR2</type>
<position>605,-145.5</position>
<input>
<ID>IN_0</ID>308 </input>
<input>
<ID>IN_1</ID>307 </input>
<output>
<ID>OUT</ID>340 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>348</ID>
<type>AI_XOR2</type>
<position>568.5,-164.5</position>
<input>
<ID>IN_0</ID>291 </input>
<input>
<ID>IN_1</ID>292 </input>
<output>
<ID>OUT</ID>296 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>349</ID>
<type>AA_LABEL</type>
<position>514.5,-151.5</position>
<gparam>LABEL_TEXT A8</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>350</ID>
<type>AA_AND2</type>
<position>554.5,-170.5</position>
<input>
<ID>IN_0</ID>285 </input>
<input>
<ID>IN_1</ID>286 </input>
<output>
<ID>OUT</ID>287 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>351</ID>
<type>AA_LABEL</type>
<position>573,-129.5</position>
<gparam>LABEL_TEXT 8-Bits Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>352</ID>
<type>DD_KEYPAD_HEX</type>
<position>522.5,-151.5</position>
<output>
<ID>OUT_0</ID>285 </output>
<output>
<ID>OUT_1</ID>291 </output>
<output>
<ID>OUT_2</ID>297 </output>
<output>
<ID>OUT_3</ID>303 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>353</ID>
<type>AE_OR2</type>
<position>582,-160.5</position>
<input>
<ID>IN_0</ID>293 </input>
<input>
<ID>IN_1</ID>294 </input>
<output>
<ID>OUT</ID>301 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>354</ID>
<type>AA_LABEL</type>
<position>514.5,-209</position>
<gparam>LABEL_TEXT B7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>355</ID>
<type>AA_AND2</type>
<position>562,-176.5</position>
<input>
<ID>IN_0</ID>290 </input>
<input>
<ID>IN_1</ID>289 </input>
<output>
<ID>OUT</ID>288 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>356</ID>
<type>AI_XOR2</type>
<position>554.5,-175.5</position>
<input>
<ID>IN_0</ID>285 </input>
<input>
<ID>IN_1</ID>286 </input>
<output>
<ID>OUT</ID>290 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>357</ID>
<type>AE_OR2</type>
<position>568,-171.5</position>
<input>
<ID>IN_0</ID>287 </input>
<input>
<ID>IN_1</ID>288 </input>
<output>
<ID>OUT</ID>295 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>358</ID>
<type>AI_XOR2</type>
<position>562,-181.5</position>
<input>
<ID>IN_0</ID>290 </input>
<input>
<ID>IN_1</ID>289 </input>
<output>
<ID>OUT</ID>337 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>359</ID>
<type>AA_AND2</type>
<position>576,-165.5</position>
<input>
<ID>IN_0</ID>296 </input>
<input>
<ID>IN_1</ID>295 </input>
<output>
<ID>OUT</ID>294 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>360</ID>
<type>DD_KEYPAD_HEX</type>
<position>522.5,-196</position>
<output>
<ID>OUT_0</ID>286 </output>
<output>
<ID>OUT_1</ID>292 </output>
<output>
<ID>OUT_2</ID>298 </output>
<output>
<ID>OUT_3</ID>304 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>361</ID>
<type>AA_AND2</type>
<position>575.5,-326.5</position>
<input>
<ID>IN_0</ID>377 </input>
<input>
<ID>IN_1</ID>376 </input>
<output>
<ID>OUT</ID>375 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>362</ID>
<type>DD_KEYPAD_HEX</type>
<position>522,-318</position>
<output>
<ID>OUT_0</ID>367 </output>
<output>
<ID>OUT_1</ID>373 </output>
<output>
<ID>OUT_2</ID>379 </output>
<output>
<ID>OUT_3</ID>385 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>363</ID>
<type>DD_KEYPAD_HEX</type>
<position>522,-273.5</position>
<output>
<ID>OUT_0</ID>366 </output>
<output>
<ID>OUT_1</ID>372 </output>
<output>
<ID>OUT_2</ID>378 </output>
<output>
<ID>OUT_3</ID>384 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<wire>
<ID>225 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>494.5,-181,494.5,-156.5</points>
<intersection>-181 1</intersection>
<intersection>-156.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>494.5,-181,500.5,-181</points>
<connection>
<GID>199</GID>
<name>IN_6</name></connection>
<intersection>494.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>470,-156.5,494.5,-156.5</points>
<connection>
<GID>181</GID>
<name>OUT</name></connection>
<intersection>494.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>397 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618,-288.5,618,-254.5</points>
<intersection>-288.5 1</intersection>
<intersection>-254.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618,-288.5,641.5,-288.5</points>
<connection>
<GID>269</GID>
<name>IN_7</name></connection>
<intersection>618 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>607.5,-254.5,618,-254.5</points>
<connection>
<GID>297</GID>
<name>OUT</name></connection>
<intersection>618 0</intersection></hsegment></shape></wire>
<wire>
<ID>396 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>617,-289.5,617,-265.5</points>
<intersection>-289.5 1</intersection>
<intersection>-265.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>617,-289.5,641.5,-289.5</points>
<connection>
<GID>269</GID>
<name>IN_6</name></connection>
<intersection>617 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>592.5,-265.5,617,-265.5</points>
<connection>
<GID>287</GID>
<name>OUT</name></connection>
<intersection>617 0</intersection></hsegment></shape></wire>
<wire>
<ID>395 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>616,-290.5,616,-279.5</points>
<intersection>-290.5 1</intersection>
<intersection>-279.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616,-290.5,641.5,-290.5</points>
<connection>
<GID>269</GID>
<name>IN_5</name></connection>
<intersection>616 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>578.5,-279.5,616,-279.5</points>
<connection>
<GID>296</GID>
<name>OUT</name></connection>
<intersection>616 0</intersection></hsegment></shape></wire>
<wire>
<ID>394 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>564.5,-291.5,641.5,-291.5</points>
<connection>
<GID>269</GID>
<name>IN_4</name></connection>
<intersection>564.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>564.5,-291.5,564.5,-290.5</points>
<connection>
<GID>307</GID>
<name>OUT</name></connection>
<intersection>-291.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>393 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>616,-306.5,616,-292.5</points>
<intersection>-306.5 2</intersection>
<intersection>-292.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616,-292.5,641.5,-292.5</points>
<connection>
<GID>269</GID>
<name>IN_3</name></connection>
<intersection>616 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>607.5,-306.5,616,-306.5</points>
<connection>
<GID>273</GID>
<name>OUT</name></connection>
<intersection>616 0</intersection></hsegment></shape></wire>
<wire>
<ID>392 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>617,-317.5,617,-293.5</points>
<intersection>-317.5 2</intersection>
<intersection>-293.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>617,-293.5,641.5,-293.5</points>
<connection>
<GID>269</GID>
<name>IN_2</name></connection>
<intersection>617 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>592.5,-317.5,617,-317.5</points>
<connection>
<GID>284</GID>
<name>OUT</name></connection>
<intersection>617 0</intersection></hsegment></shape></wire>
<wire>
<ID>391 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618,-331.5,618,-294.5</points>
<intersection>-331.5 2</intersection>
<intersection>-294.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618,-294.5,641.5,-294.5</points>
<connection>
<GID>269</GID>
<name>IN_1</name></connection>
<intersection>618 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>578.5,-331.5,618,-331.5</points>
<connection>
<GID>274</GID>
<name>OUT</name></connection>
<intersection>618 0</intersection></hsegment></shape></wire>
<wire>
<ID>390 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>619,-342.5,619,-295.5</points>
<intersection>-342.5 2</intersection>
<intersection>-295.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>619,-295.5,641.5,-295.5</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>619 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>564.5,-342.5,619,-342.5</points>
<connection>
<GID>264</GID>
<name>OUT</name></connection>
<intersection>619 0</intersection></hsegment></shape></wire>
<wire>
<ID>389 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>600,-305.5,600,-300.5</points>
<connection>
<GID>277</GID>
<name>OUT</name></connection>
<intersection>-305.5 23</intersection>
<intersection>-300.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>600,-300.5,601.5,-300.5</points>
<connection>
<GID>283</GID>
<name>IN_0</name></connection>
<intersection>600 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>600,-305.5,601.5,-305.5</points>
<connection>
<GID>273</GID>
<name>IN_0</name></connection>
<intersection>600 0</intersection></hsegment></shape></wire>
<wire>
<ID>388 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>598.5,-307.5,601.5,-307.5</points>
<connection>
<GID>273</GID>
<name>IN_1</name></connection>
<connection>
<GID>280</GID>
<name>OUT</name></connection>
<intersection>599.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>599.5,-307.5,599.5,-302.5</points>
<intersection>-307.5 1</intersection>
<intersection>-302.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>599.5,-302.5,601.5,-302.5</points>
<connection>
<GID>283</GID>
<name>IN_1</name></connection>
<intersection>599.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>387 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>607.5,-301.5,607.5,-297.5</points>
<connection>
<GID>282</GID>
<name>IN_1</name></connection>
<connection>
<GID>283</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>386 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600,-295.5,607.5,-295.5</points>
<connection>
<GID>276</GID>
<name>OUT</name></connection>
<connection>
<GID>282</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>385 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-301.5,592.5,-296.5</points>
<intersection>-301.5 2</intersection>
<intersection>-296.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>543,-301.5,594,-301.5</points>
<connection>
<GID>277</GID>
<name>IN_1</name></connection>
<intersection>543 8</intersection>
<intersection>592.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>543,-315,543,-301.5</points>
<intersection>-315 9</intersection>
<intersection>-301.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>527,-315,543,-315</points>
<connection>
<GID>362</GID>
<name>OUT_3</name></connection>
<intersection>543 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>592.5,-296.5,594,-296.5</points>
<connection>
<GID>276</GID>
<name>IN_1</name></connection>
<intersection>592.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>384 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>591,-294.5,594,-294.5</points>
<connection>
<GID>276</GID>
<name>IN_0</name></connection>
<intersection>591 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>591,-299.5,591,-294.5</points>
<intersection>-299.5 4</intersection>
<intersection>-294.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>542.5,-299.5,594,-299.5</points>
<connection>
<GID>277</GID>
<name>IN_0</name></connection>
<intersection>542.5 9</intersection>
<intersection>591 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>542.5,-299.5,542.5,-270.5</points>
<intersection>-299.5 4</intersection>
<intersection>-270.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>527,-270.5,542.5,-270.5</points>
<connection>
<GID>363</GID>
<name>OUT_3</name></connection>
<intersection>542.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>383 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585.5,-316.5,585.5,-311.5</points>
<intersection>-316.5 23</intersection>
<intersection>-311.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>585,-311.5,586.5,-311.5</points>
<connection>
<GID>279</GID>
<name>IN_0</name></connection>
<connection>
<GID>285</GID>
<name>OUT</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>585.5,-316.5,586.5,-316.5</points>
<connection>
<GID>284</GID>
<name>IN_0</name></connection>
<intersection>585.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>382 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>584.5,-318.5,586.5,-318.5</points>
<connection>
<GID>284</GID>
<name>IN_1</name></connection>
<intersection>584.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>584.5,-321.5,584.5,-313.5</points>
<connection>
<GID>268</GID>
<name>OUT</name></connection>
<intersection>-318.5 1</intersection>
<intersection>-313.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>584.5,-313.5,586.5,-313.5</points>
<connection>
<GID>279</GID>
<name>IN_1</name></connection>
<intersection>584.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>381 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-312.5,592.5,-308.5</points>
<connection>
<GID>279</GID>
<name>OUT</name></connection>
<connection>
<GID>280</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>380 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-306.5,592.5,-306.5</points>
<connection>
<GID>278</GID>
<name>OUT</name></connection>
<connection>
<GID>280</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>379 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>577,-307.5,579,-307.5</points>
<connection>
<GID>278</GID>
<name>IN_1</name></connection>
<intersection>577 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>577,-312.5,577,-307.5</points>
<intersection>-312.5 15</intersection>
<intersection>-307.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>544,-312.5,579,-312.5</points>
<connection>
<GID>285</GID>
<name>IN_1</name></connection>
<intersection>544 17</intersection>
<intersection>577 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>544,-317,544,-312.5</points>
<intersection>-317 18</intersection>
<intersection>-312.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>527,-317,544,-317</points>
<connection>
<GID>362</GID>
<name>OUT_2</name></connection>
<intersection>544 17</intersection></hsegment></shape></wire>
<wire>
<ID>378 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>544,-305.5,579,-305.5</points>
<connection>
<GID>278</GID>
<name>IN_0</name></connection>
<intersection>544 20</intersection>
<intersection>575 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>575,-310.5,575,-305.5</points>
<intersection>-310.5 16</intersection>
<intersection>-305.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>575,-310.5,579,-310.5</points>
<connection>
<GID>285</GID>
<name>IN_0</name></connection>
<intersection>575 12</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>544,-305.5,544,-272.5</points>
<intersection>-305.5 1</intersection>
<intersection>-272.5 27</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>527,-272.5,544,-272.5</points>
<connection>
<GID>363</GID>
<name>OUT_2</name></connection>
<intersection>544 20</intersection></hsegment></shape></wire>
<wire>
<ID>377 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,-330.5,571.5,-325.5</points>
<intersection>-330.5 23</intersection>
<intersection>-325.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>571,-325.5,572.5,-325.5</points>
<connection>
<GID>361</GID>
<name>IN_0</name></connection>
<connection>
<GID>272</GID>
<name>OUT</name></connection>
<intersection>571.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>571.5,-330.5,572.5,-330.5</points>
<connection>
<GID>274</GID>
<name>IN_0</name></connection>
<intersection>571.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>376 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>570.5,-332.5,572.5,-332.5</points>
<connection>
<GID>265</GID>
<name>OUT</name></connection>
<connection>
<GID>274</GID>
<name>IN_1</name></connection>
<intersection>571 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>571,-332.5,571,-327.5</points>
<intersection>-332.5 1</intersection>
<intersection>-327.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>571,-327.5,572.5,-327.5</points>
<connection>
<GID>361</GID>
<name>IN_1</name></connection>
<intersection>571 3</intersection></hsegment></shape></wire>
<wire>
<ID>375 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>578.5,-326.5,578.5,-322.5</points>
<connection>
<GID>361</GID>
<name>OUT</name></connection>
<connection>
<GID>268</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>374 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>571,-320.5,578.5,-320.5</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<connection>
<GID>281</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>373 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>563,-326.5,563,-321.5</points>
<intersection>-326.5 2</intersection>
<intersection>-321.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>544.5,-326.5,565,-326.5</points>
<connection>
<GID>272</GID>
<name>IN_1</name></connection>
<intersection>544.5 8</intersection>
<intersection>563 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>563,-321.5,565,-321.5</points>
<connection>
<GID>281</GID>
<name>IN_1</name></connection>
<intersection>563 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>544.5,-326.5,544.5,-319</points>
<intersection>-326.5 2</intersection>
<intersection>-319 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>527,-319,544.5,-319</points>
<connection>
<GID>362</GID>
<name>OUT_1</name></connection>
<intersection>544.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>372 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>545,-319.5,565,-319.5</points>
<connection>
<GID>281</GID>
<name>IN_0</name></connection>
<intersection>545 6</intersection>
<intersection>562 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>562,-324.5,562,-319.5</points>
<intersection>-324.5 4</intersection>
<intersection>-319.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>562,-324.5,565,-324.5</points>
<connection>
<GID>272</GID>
<name>IN_0</name></connection>
<intersection>562 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>545,-319.5,545,-274.5</points>
<intersection>-319.5 1</intersection>
<intersection>-274.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>527,-274.5,545,-274.5</points>
<connection>
<GID>363</GID>
<name>OUT_1</name></connection>
<intersection>545 6</intersection></hsegment></shape></wire>
<wire>
<ID>57 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,-179,269,-137.5</points>
<intersection>-179 1</intersection>
<intersection>-137.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269,-179,291.5,-179</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>263.5,-137.5,269,-137.5</points>
<connection>
<GID>22</GID>
<name>OUT</name></connection>
<intersection>269 0</intersection></hsegment></shape></wire>
<wire>
<ID>314 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>557.5,-232.5,557.5,-227.5</points>
<connection>
<GID>318</GID>
<name>OUT</name></connection>
<intersection>-232.5 23</intersection>
<intersection>-227.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>557.5,-227.5,559,-227.5</points>
<connection>
<GID>319</GID>
<name>IN_0</name></connection>
<intersection>557.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>557.5,-232.5,559,-232.5</points>
<connection>
<GID>316</GID>
<name>IN_0</name></connection>
<intersection>557.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>25 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196.5,-223.5,201,-223.5</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>196.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>196.5,-228.5,196.5,-169.5</points>
<intersection>-228.5 16</intersection>
<intersection>-223.5 1</intersection>
<intersection>-169.5 24</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>196.5,-228.5,201,-228.5</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>196.5 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>177,-169.5,196.5,-169.5</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>196.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>282 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>494,-289.5,494,-265.5</points>
<intersection>-289.5 1</intersection>
<intersection>-265.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>494,-289.5,498.5,-289.5</points>
<connection>
<GID>252</GID>
<name>IN_6</name></connection>
<intersection>494 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>469.5,-265.5,494,-265.5</points>
<connection>
<GID>234</GID>
<name>OUT</name></connection>
<intersection>494 0</intersection></hsegment></shape></wire>
<wire>
<ID>31 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>195,-212.5,215,-212.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>195 6</intersection>
<intersection>212 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>212,-217.5,212,-212.5</points>
<intersection>-217.5 4</intersection>
<intersection>-212.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>212,-217.5,215,-217.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>212 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>195,-212.5,195,-167.5</points>
<intersection>-212.5 1</intersection>
<intersection>-167.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>177,-167.5,195,-167.5</points>
<connection>
<GID>50</GID>
<name>OUT_1</name></connection>
<intersection>195 6</intersection></hsegment></shape></wire>
<wire>
<ID>288 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>565,-176.5,565,-172.5</points>
<connection>
<GID>357</GID>
<name>IN_1</name></connection>
<connection>
<GID>355</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>37 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>194,-198.5,229,-198.5</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>194 20</intersection>
<intersection>225 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>225,-203.5,225,-198.5</points>
<intersection>-203.5 16</intersection>
<intersection>-198.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>225,-203.5,229,-203.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>225 12</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>194,-198.5,194,-165.5</points>
<intersection>-198.5 1</intersection>
<intersection>-165.5 27</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>177,-165.5,194,-165.5</points>
<connection>
<GID>50</GID>
<name>OUT_2</name></connection>
<intersection>194 20</intersection></hsegment></shape></wire>
<wire>
<ID>294 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>579,-165.5,579,-161.5</points>
<connection>
<GID>359</GID>
<name>OUT</name></connection>
<connection>
<GID>353</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>43 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>241,-187.5,244,-187.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>241 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241,-192.5,241,-187.5</points>
<intersection>-192.5 4</intersection>
<intersection>-187.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>192.5,-192.5,244,-192.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>192.5 9</intersection>
<intersection>241 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>192.5,-192.5,192.5,-163.5</points>
<intersection>-192.5 4</intersection>
<intersection>-163.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>177,-163.5,192.5,-163.5</points>
<connection>
<GID>50</GID>
<name>OUT_3</name></connection>
<intersection>192.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>300 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>593,-151.5,593,-147.5</points>
<connection>
<GID>342</GID>
<name>OUT</name></connection>
<connection>
<GID>341</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>26 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>195.5,-225.5,201,-225.5</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>195.5 4</intersection>
<intersection>198.5 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>195.5,-225.5,195.5,-214</points>
<intersection>-225.5 2</intersection>
<intersection>-214 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>198.5,-230.5,198.5,-225.5</points>
<intersection>-230.5 15</intersection>
<intersection>-225.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>177,-214,195.5,-214</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>195.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>198.5,-230.5,201,-230.5</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>198.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>283 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>484.5,-288.5,498.5,-288.5</points>
<connection>
<GID>252</GID>
<name>IN_7</name></connection>
<intersection>484.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>484.5,-288.5,484.5,-254.5</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<intersection>-288.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>32 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-219.5,213,-214.5</points>
<intersection>-219.5 2</intersection>
<intersection>-214.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-219.5,215,-219.5</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>194.5 8</intersection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>213,-214.5,215,-214.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>213 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>194.5,-219.5,194.5,-212</points>
<intersection>-219.5 2</intersection>
<intersection>-212 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>177,-212,194.5,-212</points>
<connection>
<GID>49</GID>
<name>OUT_1</name></connection>
<intersection>194.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>289 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>555.5,-182.5,615.5,-182.5</points>
<connection>
<GID>358</GID>
<name>IN_1</name></connection>
<intersection>555.5 12</intersection>
<intersection>615.5 15</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>555.5,-182.5,555.5,-177.5</points>
<intersection>-182.5 1</intersection>
<intersection>-177.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>555.5,-177.5,559,-177.5</points>
<connection>
<GID>355</GID>
<name>IN_1</name></connection>
<intersection>555.5 12</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>615.5,-187.5,615.5,-182.5</points>
<intersection>-187.5 32</intersection>
<intersection>-182.5 1</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>614,-187.5,615.5,-187.5</points>
<connection>
<GID>332</GID>
<name>OUT</name></connection>
<intersection>615.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>38 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>227,-200.5,229,-200.5</points>
<connection>
<GID>33</GID>
<name>IN_1</name></connection>
<intersection>227 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>227,-205.5,227,-200.5</points>
<intersection>-205.5 15</intersection>
<intersection>-200.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>194,-205.5,229,-205.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<intersection>194 17</intersection>
<intersection>227 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>194,-210,194,-205.5</points>
<intersection>-210 18</intersection>
<intersection>-205.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>177,-210,194,-210</points>
<connection>
<GID>49</GID>
<name>OUT_2</name></connection>
<intersection>194 17</intersection></hsegment></shape></wire>
<wire>
<ID>295 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>571,-171.5,573,-171.5</points>
<connection>
<GID>346</GID>
<name>IN_1</name></connection>
<intersection>571 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>571,-171.5,571,-166.5</points>
<connection>
<GID>357</GID>
<name>OUT</name></connection>
<intersection>-171.5 1</intersection>
<intersection>-166.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>571,-166.5,573,-166.5</points>
<connection>
<GID>359</GID>
<name>IN_1</name></connection>
<intersection>571 3</intersection></hsegment></shape></wire>
<wire>
<ID>44 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242.5,-194.5,242.5,-189.5</points>
<intersection>-194.5 2</intersection>
<intersection>-189.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>193,-194.5,244,-194.5</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>193 8</intersection>
<intersection>242.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>193,-208,193,-194.5</points>
<intersection>-208 9</intersection>
<intersection>-194.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>177,-208,193,-208</points>
<connection>
<GID>49</GID>
<name>OUT_3</name></connection>
<intersection>193 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>242.5,-189.5,244,-189.5</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>242.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>301 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-157.5,587,-157.5</points>
<connection>
<GID>337</GID>
<name>IN_1</name></connection>
<intersection>585 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>585,-160.5,585,-152.5</points>
<connection>
<GID>353</GID>
<name>OUT</name></connection>
<intersection>-157.5 1</intersection>
<intersection>-152.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>585,-152.5,587,-152.5</points>
<connection>
<GID>342</GID>
<name>IN_1</name></connection>
<intersection>585 12</intersection></hsegment></shape></wire>
<wire>
<ID>36 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221.5,-223.5,221.5,-218.5</points>
<intersection>-223.5 23</intersection>
<intersection>-218.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>221,-218.5,222.5,-218.5</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>221.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>221.5,-223.5,222.5,-223.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>221.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>293 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>571.5,-159.5,579,-159.5</points>
<connection>
<GID>353</GID>
<name>IN_0</name></connection>
<connection>
<GID>340</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>35 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220.5,-225.5,222.5,-225.5</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<connection>
<GID>46</GID>
<name>OUT</name></connection>
<intersection>222 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>222,-225.5,222,-220.5</points>
<intersection>-225.5 1</intersection>
<intersection>-220.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>222,-220.5,222.5,-220.5</points>
<connection>
<GID>48</GID>
<name>IN_1</name></connection>
<intersection>222 3</intersection></hsegment></shape></wire>
<wire>
<ID>292 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>563.5,-165.5,563.5,-160.5</points>
<intersection>-165.5 2</intersection>
<intersection>-160.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>545,-165.5,565.5,-165.5</points>
<connection>
<GID>348</GID>
<name>IN_1</name></connection>
<intersection>545 8</intersection>
<intersection>563.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>563.5,-160.5,565.5,-160.5</points>
<connection>
<GID>340</GID>
<name>IN_1</name></connection>
<intersection>563.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>545,-197,545,-165.5</points>
<intersection>-197 9</intersection>
<intersection>-165.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>527.5,-197,545,-197</points>
<connection>
<GID>360</GID>
<name>OUT_1</name></connection>
<intersection>545 8</intersection></hsegment></shape></wire>
<wire>
<ID>34 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-219.5,228.5,-215.5</points>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<connection>
<GID>48</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>291 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>527.5,-152.5,565.5,-152.5</points>
<connection>
<GID>352</GID>
<name>OUT_1</name></connection>
<intersection>565.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>565.5,-163.5,565.5,-152.5</points>
<connection>
<GID>348</GID>
<name>IN_0</name></connection>
<connection>
<GID>340</GID>
<name>IN_0</name></connection>
<intersection>-152.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>30 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-234.5,207,-229.5</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<intersection>-234.5 23</intersection>
<intersection>-229.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>207,-229.5,208.5,-229.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>207,-234.5,208.5,-234.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>287 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>557.5,-170.5,565,-170.5</points>
<connection>
<GID>357</GID>
<name>IN_0</name></connection>
<connection>
<GID>350</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>29 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-236.5,208.5,-236.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>205 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>205,-236.5,205,-231.5</points>
<intersection>-236.5 1</intersection>
<intersection>-231.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>205,-231.5,208.5,-231.5</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>205 12</intersection></hsegment></shape></wire>
<wire>
<ID>286 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>546,-171.5,551.5,-171.5</points>
<connection>
<GID>350</GID>
<name>IN_1</name></connection>
<intersection>546 4</intersection>
<intersection>549 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>546,-199,546,-171.5</points>
<intersection>-199 14</intersection>
<intersection>-171.5 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>549,-176.5,549,-171.5</points>
<intersection>-176.5 15</intersection>
<intersection>-171.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>527.5,-199,546,-199</points>
<connection>
<GID>360</GID>
<name>OUT_0</name></connection>
<intersection>546 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>549,-176.5,551.5,-176.5</points>
<connection>
<GID>356</GID>
<name>IN_1</name></connection>
<intersection>549 11</intersection></hsegment></shape></wire>
<wire>
<ID>49 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>269,-235.5,269,-188.5</points>
<intersection>-235.5 2</intersection>
<intersection>-188.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>269,-188.5,291.5,-188.5</points>
<connection>
<GID>42</GID>
<name>IN_0</name></connection>
<intersection>269 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>214.5,-235.5,269,-235.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>269 0</intersection></hsegment></shape></wire>
<wire>
<ID>306 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>608,-140.5,608,-136.5</points>
<connection>
<GID>339</GID>
<name>IN_1</name></connection>
<connection>
<GID>338</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>27 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>207,-224.5,214.5,-224.5</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>28 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-230.5,214.5,-226.5</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<connection>
<GID>46</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>285 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>547,-169.5,551.5,-169.5</points>
<connection>
<GID>350</GID>
<name>IN_0</name></connection>
<intersection>547 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>547,-174.5,547,-154.5</points>
<intersection>-174.5 16</intersection>
<intersection>-169.5 1</intersection>
<intersection>-154.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>527.5,-154.5,547,-154.5</points>
<connection>
<GID>352</GID>
<name>OUT_0</name></connection>
<intersection>547 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>547,-174.5,551.5,-174.5</points>
<connection>
<GID>356</GID>
<name>IN_0</name></connection>
<intersection>547 7</intersection></hsegment></shape></wire>
<wire>
<ID>33 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221,-213.5,228.5,-213.5</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<connection>
<GID>43</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>290 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>557.5,-180.5,557.5,-175.5</points>
<connection>
<GID>356</GID>
<name>OUT</name></connection>
<intersection>-180.5 23</intersection>
<intersection>-175.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>557.5,-175.5,559,-175.5</points>
<connection>
<GID>355</GID>
<name>IN_0</name></connection>
<intersection>557.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>557.5,-180.5,559,-180.5</points>
<connection>
<GID>358</GID>
<name>IN_0</name></connection>
<intersection>557.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234.5,-211.5,236.5,-211.5</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>234.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>234.5,-214.5,234.5,-206.5</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>-211.5 1</intersection>
<intersection>-206.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>234.5,-206.5,236.5,-206.5</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>234.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>298 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>577.5,-146.5,579.5,-146.5</points>
<connection>
<GID>343</GID>
<name>IN_1</name></connection>
<intersection>577.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>577.5,-151.5,577.5,-146.5</points>
<intersection>-151.5 15</intersection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>544,-151.5,579.5,-151.5</points>
<connection>
<GID>336</GID>
<name>IN_1</name></connection>
<intersection>544 17</intersection>
<intersection>577.5 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>544,-195,544,-151.5</points>
<intersection>-195 18</intersection>
<intersection>-151.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>527.5,-195,544,-195</points>
<connection>
<GID>360</GID>
<name>OUT_2</name></connection>
<intersection>544 17</intersection></hsegment></shape></wire>
<wire>
<ID>50 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268,-224.5,268,-187.5</points>
<intersection>-224.5 2</intersection>
<intersection>-187.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268,-187.5,291.5,-187.5</points>
<connection>
<GID>42</GID>
<name>IN_1</name></connection>
<intersection>268 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228.5,-224.5,268,-224.5</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>268 0</intersection></hsegment></shape></wire>
<wire>
<ID>307 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>599,-146.5,602,-146.5</points>
<connection>
<GID>347</GID>
<name>IN_1</name></connection>
<connection>
<GID>341</GID>
<name>OUT</name></connection>
<intersection>600.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>600.5,-146.5,600.5,-141.5</points>
<intersection>-146.5 1</intersection>
<intersection>-141.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>600.5,-141.5,602,-141.5</points>
<connection>
<GID>338</GID>
<name>IN_1</name></connection>
<intersection>600.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>51 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267,-210.5,267,-186.5</points>
<intersection>-210.5 2</intersection>
<intersection>-186.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267,-186.5,291.5,-186.5</points>
<connection>
<GID>42</GID>
<name>IN_2</name></connection>
<intersection>267 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242.5,-210.5,267,-210.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>267 0</intersection></hsegment></shape></wire>
<wire>
<ID>308 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>600.5,-144.5,600.5,-139.5</points>
<connection>
<GID>344</GID>
<name>OUT</name></connection>
<intersection>-144.5 23</intersection>
<intersection>-139.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>600.5,-139.5,602,-139.5</points>
<connection>
<GID>338</GID>
<name>IN_0</name></connection>
<intersection>600.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>600.5,-144.5,602,-144.5</points>
<connection>
<GID>347</GID>
<name>IN_0</name></connection>
<intersection>600.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266,-199.5,266,-185.5</points>
<intersection>-199.5 2</intersection>
<intersection>-185.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-185.5,291.5,-185.5</points>
<connection>
<GID>42</GID>
<name>IN_3</name></connection>
<intersection>266 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>257.5,-199.5,266,-199.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>266 0</intersection></hsegment></shape></wire>
<wire>
<ID>309 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>547,-221.5,551.5,-221.5</points>
<connection>
<GID>322</GID>
<name>IN_0</name></connection>
<intersection>547 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>547,-226.5,547,-167.5</points>
<intersection>-226.5 16</intersection>
<intersection>-221.5 1</intersection>
<intersection>-167.5 24</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>547,-226.5,551.5,-226.5</points>
<connection>
<GID>318</GID>
<name>IN_0</name></connection>
<intersection>547 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>527.5,-167.5,547,-167.5</points>
<connection>
<GID>313</GID>
<name>OUT_0</name></connection>
<intersection>547 7</intersection></hsegment></shape></wire>
<wire>
<ID>53 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>214.5,-184.5,291.5,-184.5</points>
<connection>
<GID>42</GID>
<name>IN_4</name></connection>
<intersection>214.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>214.5,-184.5,214.5,-183.5</points>
<connection>
<GID>3</GID>
<name>OUT</name></connection>
<intersection>-184.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>310 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>546,-223.5,551.5,-223.5</points>
<connection>
<GID>322</GID>
<name>IN_1</name></connection>
<intersection>546 4</intersection>
<intersection>549 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>546,-223.5,546,-212</points>
<intersection>-223.5 2</intersection>
<intersection>-212 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>549,-228.5,549,-223.5</points>
<intersection>-228.5 15</intersection>
<intersection>-223.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>527.5,-212,546,-212</points>
<connection>
<GID>314</GID>
<name>OUT_0</name></connection>
<intersection>546 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>549,-228.5,551.5,-228.5</points>
<connection>
<GID>318</GID>
<name>IN_1</name></connection>
<intersection>549 11</intersection></hsegment></shape></wire>
<wire>
<ID>54 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266,-183.5,266,-172.5</points>
<intersection>-183.5 1</intersection>
<intersection>-172.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>266,-183.5,291.5,-183.5</points>
<connection>
<GID>42</GID>
<name>IN_5</name></connection>
<intersection>266 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>228.5,-172.5,266,-172.5</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>266 0</intersection></hsegment></shape></wire>
<wire>
<ID>311 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>557.5,-222.5,565,-222.5</points>
<connection>
<GID>322</GID>
<name>OUT</name></connection>
<connection>
<GID>317</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>55 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>267,-182.5,267,-158.5</points>
<intersection>-182.5 1</intersection>
<intersection>-158.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>267,-182.5,291.5,-182.5</points>
<connection>
<GID>42</GID>
<name>IN_6</name></connection>
<intersection>267 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>242.5,-158.5,267,-158.5</points>
<connection>
<GID>24</GID>
<name>OUT</name></connection>
<intersection>267 0</intersection></hsegment></shape></wire>
<wire>
<ID>312 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>565,-228.5,565,-224.5</points>
<connection>
<GID>319</GID>
<name>OUT</name></connection>
<connection>
<GID>317</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>56 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>268,-181.5,268,-147.5</points>
<intersection>-181.5 1</intersection>
<intersection>-147.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>268,-181.5,291.5,-181.5</points>
<connection>
<GID>42</GID>
<name>IN_7</name></connection>
<intersection>268 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>257.5,-147.5,268,-147.5</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>268 0</intersection></hsegment></shape></wire>
<wire>
<ID>313 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>555.5,-236.5,613.5,-236.5</points>
<intersection>555.5 12</intersection>
<intersection>559 19</intersection>
<intersection>613.5 17</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>555.5,-236.5,555.5,-229.5</points>
<intersection>-236.5 1</intersection>
<intersection>-229.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>555.5,-229.5,559,-229.5</points>
<connection>
<GID>319</GID>
<name>IN_1</name></connection>
<intersection>555.5 12</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>613.5,-244.5,613.5,-236.5</points>
<connection>
<GID>289</GID>
<name>OUT</name></connection>
<intersection>-236.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>559,-236.5,559,-234.5</points>
<connection>
<GID>316</GID>
<name>IN_1</name></connection>
<intersection>-236.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>48 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-198.5,250,-193.5</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>-198.5 23</intersection>
<intersection>-193.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>250,-193.5,251.5,-193.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>250,-198.5,251.5,-198.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>250 0</intersection></hsegment></shape></wire>
<wire>
<ID>305 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600.5,-134.5,608,-134.5</points>
<connection>
<GID>345</GID>
<name>OUT</name></connection>
<connection>
<GID>339</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>47 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>248.5,-200.5,251.5,-200.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>248.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>248.5,-200.5,248.5,-195.5</points>
<intersection>-200.5 1</intersection>
<intersection>-195.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>248.5,-195.5,251.5,-195.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>248.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>304 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>593,-140.5,593,-135.5</points>
<intersection>-140.5 2</intersection>
<intersection>-135.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>543.5,-140.5,594.5,-140.5</points>
<connection>
<GID>344</GID>
<name>IN_1</name></connection>
<intersection>543.5 8</intersection>
<intersection>593 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>543.5,-193,543.5,-140.5</points>
<intersection>-193 9</intersection>
<intersection>-140.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>527.5,-193,543.5,-193</points>
<connection>
<GID>360</GID>
<name>OUT_3</name></connection>
<intersection>543.5 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>593,-135.5,594.5,-135.5</points>
<connection>
<GID>345</GID>
<name>IN_1</name></connection>
<intersection>593 0</intersection></hsegment></shape></wire>
<wire>
<ID>45 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>250,-188.5,257.5,-188.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<connection>
<GID>35</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>302 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585.5,-155.5,585.5,-150.5</points>
<connection>
<GID>336</GID>
<name>OUT</name></connection>
<intersection>-155.5 23</intersection>
<intersection>-150.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>585.5,-150.5,587,-150.5</points>
<connection>
<GID>342</GID>
<name>IN_0</name></connection>
<intersection>585.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>585.5,-155.5,587,-155.5</points>
<connection>
<GID>337</GID>
<name>IN_0</name></connection>
<intersection>585.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235,-199.5,242.5,-199.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<connection>
<GID>33</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>296 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571.5,-169.5,571.5,-164.5</points>
<connection>
<GID>348</GID>
<name>OUT</name></connection>
<intersection>-169.5 23</intersection>
<intersection>-164.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>571.5,-164.5,573,-164.5</points>
<connection>
<GID>359</GID>
<name>IN_0</name></connection>
<intersection>571.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>571.5,-169.5,573,-169.5</points>
<connection>
<GID>346</GID>
<name>IN_0</name></connection>
<intersection>571.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>42 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235.5,-209.5,235.5,-204.5</points>
<intersection>-209.5 23</intersection>
<intersection>-204.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>235,-204.5,236.5,-204.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>235.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>235.5,-209.5,236.5,-209.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>235.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>299 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585.5,-145.5,593,-145.5</points>
<connection>
<GID>343</GID>
<name>OUT</name></connection>
<connection>
<GID>341</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>40 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242.5,-205.5,242.5,-201.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<connection>
<GID>32</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>297 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>527.5,-150.5,579.5,-150.5</points>
<connection>
<GID>352</GID>
<name>OUT_2</name></connection>
<intersection>574.5 20</intersection>
<intersection>579.5 23</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>574.5,-150.5,574.5,-144.5</points>
<intersection>-150.5 1</intersection>
<intersection>-144.5 22</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>574.5,-144.5,579.5,-144.5</points>
<connection>
<GID>343</GID>
<name>IN_0</name></connection>
<intersection>574.5 20</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>579.5,-150.5,579.5,-149.5</points>
<connection>
<GID>336</GID>
<name>IN_0</name></connection>
<intersection>-150.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>46 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257.5,-194.5,257.5,-190.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<connection>
<GID>29</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>303 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>543,-133.5,594.5,-133.5</points>
<connection>
<GID>345</GID>
<name>IN_0</name></connection>
<intersection>543 6</intersection>
<intersection>592 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>592,-138.5,592,-133.5</points>
<intersection>-138.5 4</intersection>
<intersection>-133.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>592,-138.5,594.5,-138.5</points>
<connection>
<GID>344</GID>
<name>IN_0</name></connection>
<intersection>592 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>543,-148.5,543,-133.5</points>
<intersection>-148.5 8</intersection>
<intersection>-133.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>527.5,-148.5,543,-148.5</points>
<connection>
<GID>352</GID>
<name>OUT_3</name></connection>
<intersection>543 6</intersection></hsegment></shape></wire>
<wire>
<ID>5 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>205,-186,265,-186</points>
<intersection>205 12</intersection>
<intersection>208.5 19</intersection>
<intersection>265 15</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>205,-186,205,-179.5</points>
<intersection>-186 1</intersection>
<intersection>-179.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>205,-179.5,208.5,-179.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>205 12</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>265,-189.5,265,-186</points>
<intersection>-189.5 32</intersection>
<intersection>-186 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>208.5,-186,208.5,-184.5</points>
<connection>
<GID>3</GID>
<name>IN_1</name></connection>
<intersection>-186 1</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>263.5,-189.5,265,-189.5</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>265 15</intersection></hsegment></shape></wire>
<wire>
<ID>262 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>447.5,-332.5,449.5,-332.5</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<connection>
<GID>247</GID>
<name>IN_1</name></connection>
<intersection>449 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>449,-332.5,449,-327.5</points>
<intersection>-332.5 1</intersection>
<intersection>-327.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>449,-327.5,449.5,-327.5</points>
<connection>
<GID>258</GID>
<name>IN_1</name></connection>
<intersection>449 3</intersection></hsegment></shape></wire>
<wire>
<ID>13 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-152.5,229,-152.5</points>
<connection>
<GID>9</GID>
<name>OUT_2</name></connection>
<intersection>224 20</intersection>
<intersection>229 23</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>224,-152.5,224,-146.5</points>
<intersection>-152.5 1</intersection>
<intersection>-146.5 22</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>224,-146.5,229,-146.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>224 20</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>229,-152.5,229,-151.5</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>-152.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>270 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>468,-294.5,471,-294.5</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>468 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>468,-299.5,468,-294.5</points>
<intersection>-299.5 4</intersection>
<intersection>-294.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>419.5,-299.5,471,-299.5</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>419.5 9</intersection>
<intersection>468 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>419.5,-299.5,419.5,-270.5</points>
<intersection>-299.5 4</intersection>
<intersection>-270.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>404,-270.5,419.5,-270.5</points>
<connection>
<GID>260</GID>
<name>OUT_3</name></connection>
<intersection>419.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>14 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>227,-148.5,229,-148.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>227 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>227,-153.5,227,-148.5</points>
<intersection>-153.5 15</intersection>
<intersection>-148.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>193.5,-153.5,229,-153.5</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>193.5 17</intersection>
<intersection>227 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>193.5,-197,193.5,-153.5</points>
<intersection>-197 18</intersection>
<intersection>-153.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>177,-197,193.5,-197</points>
<connection>
<GID>1</GID>
<name>OUT_2</name></connection>
<intersection>193.5 17</intersection></hsegment></shape></wire>
<wire>
<ID>271 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>469.5,-301.5,469.5,-296.5</points>
<intersection>-301.5 2</intersection>
<intersection>-296.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>420,-301.5,471,-301.5</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>420 8</intersection>
<intersection>469.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>420,-315,420,-301.5</points>
<intersection>-315 9</intersection>
<intersection>-301.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>404,-315,420,-315</points>
<connection>
<GID>259</GID>
<name>OUT_3</name></connection>
<intersection>420 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>469.5,-296.5,471,-296.5</points>
<connection>
<GID>245</GID>
<name>IN_1</name></connection>
<intersection>469.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>235,-157.5,235,-152.5</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<intersection>-157.5 23</intersection>
<intersection>-152.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>235,-152.5,236.5,-152.5</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>235,-157.5,236.5,-157.5</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>235 0</intersection></hsegment></shape></wire>
<wire>
<ID>275 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>477,-305.5,477,-300.5</points>
<connection>
<GID>244</GID>
<name>OUT</name></connection>
<intersection>-305.5 23</intersection>
<intersection>-300.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>477,-300.5,478.5,-300.5</points>
<connection>
<GID>238</GID>
<name>IN_0</name></connection>
<intersection>477 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>477,-305.5,478.5,-305.5</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>477 0</intersection></hsegment></shape></wire>
<wire>
<ID>17 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>234.5,-159.5,236.5,-159.5</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>234.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>234.5,-162.5,234.5,-154.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>-159.5 1</intersection>
<intersection>-154.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>234.5,-154.5,236.5,-154.5</points>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>234.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>274 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>475.5,-307.5,478.5,-307.5</points>
<connection>
<GID>241</GID>
<name>OUT</name></connection>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<intersection>476.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>476.5,-307.5,476.5,-302.5</points>
<intersection>-307.5 1</intersection>
<intersection>-302.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>476.5,-302.5,478.5,-302.5</points>
<connection>
<GID>238</GID>
<name>IN_1</name></connection>
<intersection>476.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>24 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>250,-146.5,250,-141.5</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>-146.5 23</intersection>
<intersection>-141.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>250,-141.5,251.5,-141.5</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>250 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>250,-146.5,251.5,-146.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>250 0</intersection></hsegment></shape></wire>
<wire>
<ID>281 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>493,-290.5,493,-279.5</points>
<intersection>-290.5 1</intersection>
<intersection>-279.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>493,-290.5,498.5,-290.5</points>
<connection>
<GID>252</GID>
<name>IN_5</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>455.5,-279.5,493,-279.5</points>
<connection>
<GID>225</GID>
<name>OUT</name></connection>
<intersection>493 0</intersection></hsegment></shape></wire>
<wire>
<ID>23 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>248.5,-148.5,251.5,-148.5</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>250 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>250,-148.5,250,-143.5</points>
<intersection>-148.5 1</intersection>
<intersection>-143.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>250,-143.5,251.5,-143.5</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>250 3</intersection></hsegment></shape></wire>
<wire>
<ID>280 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>441.5,-291.5,498.5,-291.5</points>
<connection>
<GID>252</GID>
<name>IN_4</name></connection>
<intersection>441.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>441.5,-291.5,441.5,-290.5</points>
<connection>
<GID>213</GID>
<name>OUT</name></connection>
<intersection>-291.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>22 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>257.5,-142.5,257.5,-138.5</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<connection>
<GID>23</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>279 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>493,-306.5,493,-292.5</points>
<intersection>-306.5 2</intersection>
<intersection>-292.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>493,-292.5,498.5,-292.5</points>
<connection>
<GID>252</GID>
<name>IN_3</name></connection>
<intersection>493 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>484.5,-306.5,493,-306.5</points>
<connection>
<GID>248</GID>
<name>OUT</name></connection>
<intersection>493 0</intersection></hsegment></shape></wire>
<wire>
<ID>21 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>250,-136.5,257.5,-136.5</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<connection>
<GID>22</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>278 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>494,-317.5,494,-293.5</points>
<intersection>-317.5 2</intersection>
<intersection>-293.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>494,-293.5,498.5,-293.5</points>
<connection>
<GID>252</GID>
<name>IN_2</name></connection>
<intersection>494 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>469.5,-317.5,494,-317.5</points>
<connection>
<GID>237</GID>
<name>OUT</name></connection>
<intersection>494 0</intersection></hsegment></shape></wire>
<wire>
<ID>7 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-154.5,215,-154.5</points>
<connection>
<GID>9</GID>
<name>OUT_1</name></connection>
<intersection>215 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>215,-165.5,215,-154.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>-154.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>264 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>421,-305.5,456,-305.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>421 20</intersection>
<intersection>452 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>452,-310.5,452,-305.5</points>
<intersection>-310.5 16</intersection>
<intersection>-305.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>452,-310.5,456,-310.5</points>
<connection>
<GID>236</GID>
<name>IN_0</name></connection>
<intersection>452 12</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>421,-305.5,421,-272.5</points>
<intersection>-305.5 1</intersection>
<intersection>-272.5 27</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>404,-272.5,421,-272.5</points>
<connection>
<GID>260</GID>
<name>OUT_2</name></connection>
<intersection>421 20</intersection></hsegment></shape></wire>
<wire>
<ID>8 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>213,-167.5,213,-162.5</points>
<intersection>-167.5 2</intersection>
<intersection>-162.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>194.5,-167.5,215,-167.5</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>194.5 8</intersection>
<intersection>213 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>213,-162.5,215,-162.5</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>213 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>194.5,-199,194.5,-167.5</points>
<intersection>-199 9</intersection>
<intersection>-167.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>177,-199,194.5,-199</points>
<connection>
<GID>1</GID>
<name>OUT_1</name></connection>
<intersection>194.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>265 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>454,-307.5,456,-307.5</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<intersection>454 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>454,-312.5,454,-307.5</points>
<intersection>-312.5 15</intersection>
<intersection>-307.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>421,-312.5,456,-312.5</points>
<connection>
<GID>236</GID>
<name>IN_1</name></connection>
<intersection>421 17</intersection>
<intersection>454 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>421,-317,421,-312.5</points>
<intersection>-317 18</intersection>
<intersection>-312.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>404,-317,421,-317</points>
<connection>
<GID>259</GID>
<name>OUT_2</name></connection>
<intersection>421 17</intersection></hsegment></shape></wire>
<wire>
<ID>9 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>221,-161.5,228.5,-161.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<connection>
<GID>21</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>266 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>462,-306.5,469.5,-306.5</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<connection>
<GID>241</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>15 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>235,-147.5,242.5,-147.5</points>
<connection>
<GID>18</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>272 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477,-295.5,484.5,-295.5</points>
<connection>
<GID>245</GID>
<name>OUT</name></connection>
<connection>
<GID>239</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>16 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242.5,-153.5,242.5,-149.5</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<connection>
<GID>20</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>273 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484.5,-301.5,484.5,-297.5</points>
<connection>
<GID>238</GID>
<name>OUT</name></connection>
<connection>
<GID>239</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>19 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>192.5,-135.5,244,-135.5</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>192.5 6</intersection>
<intersection>241.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>241.5,-140.5,241.5,-135.5</points>
<intersection>-140.5 4</intersection>
<intersection>-135.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>241.5,-140.5,244,-140.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>241.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>192.5,-150.5,192.5,-135.5</points>
<intersection>-150.5 8</intersection>
<intersection>-135.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>177,-150.5,192.5,-150.5</points>
<connection>
<GID>9</GID>
<name>OUT_3</name></connection>
<intersection>192.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>276 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>496,-342.5,496,-295.5</points>
<intersection>-342.5 2</intersection>
<intersection>-295.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>496,-295.5,498.5,-295.5</points>
<connection>
<GID>252</GID>
<name>IN_0</name></connection>
<intersection>496 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>441.5,-342.5,496,-342.5</points>
<connection>
<GID>257</GID>
<name>OUT</name></connection>
<intersection>496 0</intersection></hsegment></shape></wire>
<wire>
<ID>20 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>242.5,-142.5,242.5,-137.5</points>
<intersection>-142.5 2</intersection>
<intersection>-137.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>193,-142.5,244,-142.5</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>193 8</intersection>
<intersection>242.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>193,-195,193,-142.5</points>
<intersection>-195 9</intersection>
<intersection>-142.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>177,-195,193,-195</points>
<connection>
<GID>1</GID>
<name>OUT_3</name></connection>
<intersection>193 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>242.5,-137.5,244,-137.5</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>242.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>277 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>495,-331.5,495,-294.5</points>
<intersection>-331.5 2</intersection>
<intersection>-294.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>495,-294.5,498.5,-294.5</points>
<connection>
<GID>252</GID>
<name>IN_1</name></connection>
<intersection>495 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>455.5,-331.5,495,-331.5</points>
<connection>
<GID>247</GID>
<name>OUT</name></connection>
<intersection>495 0</intersection></hsegment></shape></wire>
<wire>
<ID>12 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>221,-171.5,221,-166.5</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>-171.5 23</intersection>
<intersection>-166.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>221,-166.5,222.5,-166.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>221 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>221,-171.5,222.5,-171.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<intersection>221 0</intersection></hsegment></shape></wire>
<wire>
<ID>269 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462.5,-316.5,462.5,-311.5</points>
<intersection>-316.5 23</intersection>
<intersection>-311.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>462,-311.5,463.5,-311.5</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<connection>
<GID>236</GID>
<name>OUT</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>462.5,-316.5,463.5,-316.5</points>
<connection>
<GID>237</GID>
<name>IN_0</name></connection>
<intersection>462.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>220.5,-173.5,222.5,-173.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<intersection>220.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>220.5,-173.5,220.5,-168.5</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>-173.5 1</intersection>
<intersection>-168.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>220.5,-168.5,222.5,-168.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>220.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>268 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>461.5,-318.5,463.5,-318.5</points>
<connection>
<GID>237</GID>
<name>IN_1</name></connection>
<intersection>461.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>461.5,-321.5,461.5,-313.5</points>
<connection>
<GID>253</GID>
<name>OUT</name></connection>
<intersection>-318.5 1</intersection>
<intersection>-313.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>461.5,-313.5,463.5,-313.5</points>
<connection>
<GID>242</GID>
<name>IN_1</name></connection>
<intersection>461.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>1 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>196.5,-171.5,201,-171.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>196.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>196.5,-176.5,196.5,-156.5</points>
<intersection>-176.5 16</intersection>
<intersection>-171.5 1</intersection>
<intersection>-156.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>177,-156.5,196.5,-156.5</points>
<connection>
<GID>9</GID>
<name>OUT_0</name></connection>
<intersection>196.5 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>196.5,-176.5,201,-176.5</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>196.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>258 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>422,-319.5,442,-319.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>422 6</intersection>
<intersection>439 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>439,-324.5,439,-319.5</points>
<intersection>-324.5 4</intersection>
<intersection>-319.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>439,-324.5,442,-324.5</points>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>439 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>422,-319.5,422,-274.5</points>
<intersection>-319.5 1</intersection>
<intersection>-274.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>404,-274.5,422,-274.5</points>
<connection>
<GID>260</GID>
<name>OUT_1</name></connection>
<intersection>422 6</intersection></hsegment></shape></wire>
<wire>
<ID>2 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>195.5,-173.5,201,-173.5</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>195.5 4</intersection>
<intersection>198.5 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>195.5,-201,195.5,-173.5</points>
<intersection>-201 14</intersection>
<intersection>-173.5 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>198.5,-178.5,198.5,-173.5</points>
<intersection>-178.5 15</intersection>
<intersection>-173.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>177,-201,195.5,-201</points>
<connection>
<GID>1</GID>
<name>OUT_0</name></connection>
<intersection>195.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>198.5,-178.5,201,-178.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>198.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>259 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>440,-326.5,440,-321.5</points>
<intersection>-326.5 2</intersection>
<intersection>-321.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>421.5,-326.5,442,-326.5</points>
<connection>
<GID>249</GID>
<name>IN_1</name></connection>
<intersection>421.5 8</intersection>
<intersection>440 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440,-321.5,442,-321.5</points>
<connection>
<GID>240</GID>
<name>IN_1</name></connection>
<intersection>440 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>421.5,-326.5,421.5,-319</points>
<intersection>-326.5 2</intersection>
<intersection>-319 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>404,-319,421.5,-319</points>
<connection>
<GID>259</GID>
<name>OUT_1</name></connection>
<intersection>421.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>3 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>207,-172.5,214.5,-172.5</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<connection>
<GID>11</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>260 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>448,-320.5,455.5,-320.5</points>
<connection>
<GID>240</GID>
<name>OUT</name></connection>
<connection>
<GID>253</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>228.5,-167.5,228.5,-163.5</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>8</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>267 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>469.5,-312.5,469.5,-308.5</points>
<connection>
<GID>241</GID>
<name>IN_1</name></connection>
<connection>
<GID>242</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>6 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>207,-182.5,207,-177.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>-182.5 23</intersection>
<intersection>-177.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>207,-177.5,208.5,-177.5</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>207,-182.5,208.5,-182.5</points>
<connection>
<GID>3</GID>
<name>IN_0</name></connection>
<intersection>207 0</intersection></hsegment></shape></wire>
<wire>
<ID>263 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448.5,-330.5,448.5,-325.5</points>
<intersection>-330.5 23</intersection>
<intersection>-325.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>448,-325.5,449.5,-325.5</points>
<connection>
<GID>249</GID>
<name>OUT</name></connection>
<connection>
<GID>258</GID>
<name>IN_0</name></connection>
<intersection>448.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>448.5,-330.5,449.5,-330.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<intersection>448.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>214.5,-178.5,214.5,-174.5</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<connection>
<GID>6</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>261 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455.5,-326.5,455.5,-322.5</points>
<connection>
<GID>258</GID>
<name>OUT</name></connection>
<connection>
<GID>253</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>171 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>424,-169.5,428.5,-169.5</points>
<connection>
<GID>168</GID>
<name>IN_0</name></connection>
<intersection>424 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>424,-174.5,424,-154.5</points>
<intersection>-174.5 16</intersection>
<intersection>-169.5 1</intersection>
<intersection>-154.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>404.5,-154.5,424,-154.5</points>
<connection>
<GID>166</GID>
<name>OUT_0</name></connection>
<intersection>424 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>424,-174.5,428.5,-174.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>424 7</intersection></hsegment></shape></wire>
<wire>
<ID>172 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>423,-171.5,428.5,-171.5</points>
<connection>
<GID>168</GID>
<name>IN_1</name></connection>
<intersection>423 4</intersection>
<intersection>426 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>423,-199,423,-171.5</points>
<intersection>-199 14</intersection>
<intersection>-171.5 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>426,-176.5,426,-171.5</points>
<intersection>-176.5 15</intersection>
<intersection>-171.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>404.5,-199,423,-199</points>
<connection>
<GID>158</GID>
<name>OUT_0</name></connection>
<intersection>423 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>426,-176.5,428.5,-176.5</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>426 11</intersection></hsegment></shape></wire>
<wire>
<ID>173 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>434.5,-170.5,442,-170.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<connection>
<GID>168</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>174 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>442,-176.5,442,-172.5</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<connection>
<GID>163</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>175 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432.5,-184,492.5,-184</points>
<intersection>432.5 12</intersection>
<intersection>436 19</intersection>
<intersection>492.5 15</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>432.5,-184,432.5,-177.5</points>
<intersection>-184 1</intersection>
<intersection>-177.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>432.5,-177.5,436,-177.5</points>
<connection>
<GID>163</GID>
<name>IN_1</name></connection>
<intersection>432.5 12</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>492.5,-187.5,492.5,-184</points>
<intersection>-187.5 32</intersection>
<intersection>-184 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>436,-184,436,-182.5</points>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>-184 1</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>491,-187.5,492.5,-187.5</points>
<connection>
<GID>186</GID>
<name>OUT</name></connection>
<intersection>492.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>176 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,-180.5,434.5,-175.5</points>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<intersection>-180.5 23</intersection>
<intersection>-175.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>434.5,-175.5,436,-175.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>434.5,-180.5,436,-180.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>434.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>177 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>404.5,-152.5,442.5,-152.5</points>
<connection>
<GID>166</GID>
<name>OUT_1</name></connection>
<intersection>442.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>442.5,-163.5,442.5,-152.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>-152.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>178 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>440.5,-165.5,440.5,-160.5</points>
<intersection>-165.5 2</intersection>
<intersection>-160.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>422,-165.5,442.5,-165.5</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>422 8</intersection>
<intersection>440.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440.5,-160.5,442.5,-160.5</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<intersection>440.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>422,-197,422,-165.5</points>
<intersection>-197 9</intersection>
<intersection>-165.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>404.5,-197,422,-197</points>
<connection>
<GID>158</GID>
<name>OUT_1</name></connection>
<intersection>422 8</intersection></hsegment></shape></wire>
<wire>
<ID>179 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>448.5,-159.5,456,-159.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>180 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,-165.5,456,-161.5</points>
<connection>
<GID>159</GID>
<name>OUT</name></connection>
<connection>
<GID>165</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>181 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>448,-171.5,450,-171.5</points>
<connection>
<GID>172</GID>
<name>IN_1</name></connection>
<intersection>448 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>448,-171.5,448,-166.5</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>-171.5 1</intersection>
<intersection>-166.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>448,-166.5,450,-166.5</points>
<connection>
<GID>159</GID>
<name>IN_1</name></connection>
<intersection>448 3</intersection></hsegment></shape></wire>
<wire>
<ID>182 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448.5,-169.5,448.5,-164.5</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<intersection>-169.5 23</intersection>
<intersection>-164.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>448.5,-164.5,450,-164.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>448.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>448.5,-169.5,450,-169.5</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>448.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>183 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>404.5,-150.5,456.5,-150.5</points>
<connection>
<GID>166</GID>
<name>OUT_2</name></connection>
<intersection>451.5 20</intersection>
<intersection>456.5 23</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>451.5,-150.5,451.5,-144.5</points>
<intersection>-150.5 1</intersection>
<intersection>-144.5 22</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>451.5,-144.5,456.5,-144.5</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>451.5 20</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>456.5,-150.5,456.5,-149.5</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<intersection>-150.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>184 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>454.5,-146.5,456.5,-146.5</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>454.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>454.5,-151.5,454.5,-146.5</points>
<intersection>-151.5 15</intersection>
<intersection>-146.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>421,-151.5,456.5,-151.5</points>
<connection>
<GID>182</GID>
<name>IN_1</name></connection>
<intersection>421 17</intersection>
<intersection>454.5 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>421,-195,421,-151.5</points>
<intersection>-195 18</intersection>
<intersection>-151.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>404.5,-195,421,-195</points>
<connection>
<GID>158</GID>
<name>OUT_2</name></connection>
<intersection>421 17</intersection></hsegment></shape></wire>
<wire>
<ID>185 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>462.5,-145.5,470,-145.5</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<connection>
<GID>177</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>186 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>470,-151.5,470,-147.5</points>
<connection>
<GID>176</GID>
<name>OUT</name></connection>
<connection>
<GID>177</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>187 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>462,-157.5,464,-157.5</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<intersection>462 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>462,-160.5,462,-152.5</points>
<connection>
<GID>165</GID>
<name>OUT</name></connection>
<intersection>-157.5 1</intersection>
<intersection>-152.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>462,-152.5,464,-152.5</points>
<connection>
<GID>176</GID>
<name>IN_1</name></connection>
<intersection>462 12</intersection></hsegment></shape></wire>
<wire>
<ID>188 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462.5,-155.5,462.5,-150.5</points>
<connection>
<GID>182</GID>
<name>OUT</name></connection>
<intersection>-155.5 23</intersection>
<intersection>-150.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>462.5,-150.5,464,-150.5</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>462.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>462.5,-155.5,464,-155.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>462.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>189 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>420,-133.5,471.5,-133.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>420 6</intersection>
<intersection>469 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>469,-138.5,469,-133.5</points>
<intersection>-138.5 4</intersection>
<intersection>-133.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>469,-138.5,471.5,-138.5</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<intersection>469 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>420,-148.5,420,-133.5</points>
<intersection>-148.5 8</intersection>
<intersection>-133.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>404.5,-148.5,420,-148.5</points>
<connection>
<GID>166</GID>
<name>OUT_3</name></connection>
<intersection>420 6</intersection></hsegment></shape></wire>
<wire>
<ID>190 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>470,-140.5,470,-135.5</points>
<intersection>-140.5 2</intersection>
<intersection>-135.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>420.5,-140.5,471.5,-140.5</points>
<connection>
<GID>174</GID>
<name>IN_1</name></connection>
<intersection>420.5 8</intersection>
<intersection>470 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>420.5,-193,420.5,-140.5</points>
<intersection>-193 9</intersection>
<intersection>-140.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>404.5,-193,420.5,-193</points>
<connection>
<GID>158</GID>
<name>OUT_3</name></connection>
<intersection>420.5 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>470,-135.5,471.5,-135.5</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>470 0</intersection></hsegment></shape></wire>
<wire>
<ID>191 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477.5,-134.5,485,-134.5</points>
<connection>
<GID>173</GID>
<name>OUT</name></connection>
<connection>
<GID>179</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>192 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>485,-140.5,485,-136.5</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<connection>
<GID>180</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>193 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>476,-146.5,479,-146.5</points>
<connection>
<GID>171</GID>
<name>IN_1</name></connection>
<connection>
<GID>177</GID>
<name>OUT</name></connection>
<intersection>477.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>477.5,-146.5,477.5,-141.5</points>
<intersection>-146.5 1</intersection>
<intersection>-141.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>477.5,-141.5,479,-141.5</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>477.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>194 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>477.5,-144.5,477.5,-139.5</points>
<connection>
<GID>174</GID>
<name>OUT</name></connection>
<intersection>-144.5 23</intersection>
<intersection>-139.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>477.5,-139.5,479,-139.5</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>477.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>477.5,-144.5,479,-144.5</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>477.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>195 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>424,-221.5,428.5,-221.5</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>424 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>424,-226.5,424,-167.5</points>
<intersection>-226.5 16</intersection>
<intersection>-221.5 1</intersection>
<intersection>-167.5 24</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>424,-226.5,428.5,-226.5</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>424 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>404.5,-167.5,424,-167.5</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<intersection>424 7</intersection></hsegment></shape></wire>
<wire>
<ID>196 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>423,-223.5,428.5,-223.5</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>423 4</intersection>
<intersection>426 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>423,-223.5,423,-212</points>
<intersection>-223.5 2</intersection>
<intersection>-212 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>426,-228.5,426,-223.5</points>
<intersection>-228.5 15</intersection>
<intersection>-223.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>404.5,-212,423,-212</points>
<connection>
<GID>206</GID>
<name>OUT_0</name></connection>
<intersection>423 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>426,-228.5,428.5,-228.5</points>
<connection>
<GID>202</GID>
<name>IN_1</name></connection>
<intersection>426 11</intersection></hsegment></shape></wire>
<wire>
<ID>197 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>434.5,-222.5,442,-222.5</points>
<connection>
<GID>197</GID>
<name>OUT</name></connection>
<connection>
<GID>203</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>198 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>442,-228.5,442,-224.5</points>
<connection>
<GID>201</GID>
<name>OUT</name></connection>
<connection>
<GID>203</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>199 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432.5,-236.5,490.5,-236.5</points>
<intersection>432.5 12</intersection>
<intersection>436 19</intersection>
<intersection>490.5 17</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>432.5,-236.5,432.5,-229.5</points>
<intersection>-236.5 1</intersection>
<intersection>-229.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>432.5,-229.5,436,-229.5</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>432.5 12</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>490.5,-244.5,490.5,-236.5</points>
<connection>
<GID>232</GID>
<name>OUT</name></connection>
<intersection>-236.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>436,-236.5,436,-234.5</points>
<connection>
<GID>204</GID>
<name>IN_1</name></connection>
<intersection>-236.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>200 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434.5,-232.5,434.5,-227.5</points>
<connection>
<GID>202</GID>
<name>OUT</name></connection>
<intersection>-232.5 23</intersection>
<intersection>-227.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>434.5,-227.5,436,-227.5</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>434.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>434.5,-232.5,436,-232.5</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>434.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>201 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>422.5,-210.5,442.5,-210.5</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>422.5 6</intersection>
<intersection>439.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>439.5,-215.5,439.5,-210.5</points>
<intersection>-215.5 4</intersection>
<intersection>-210.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>439.5,-215.5,442.5,-215.5</points>
<connection>
<GID>196</GID>
<name>IN_0</name></connection>
<intersection>439.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>422.5,-210.5,422.5,-165.5</points>
<intersection>-210.5 1</intersection>
<intersection>-165.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>404.5,-165.5,422.5,-165.5</points>
<connection>
<GID>207</GID>
<name>OUT_1</name></connection>
<intersection>422.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>202 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>440.5,-217.5,440.5,-212.5</points>
<intersection>-217.5 2</intersection>
<intersection>-212.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>422,-217.5,442.5,-217.5</points>
<connection>
<GID>196</GID>
<name>IN_1</name></connection>
<intersection>422 8</intersection>
<intersection>440.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440.5,-212.5,442.5,-212.5</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>440.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>422,-217.5,422,-210</points>
<intersection>-217.5 2</intersection>
<intersection>-210 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>404.5,-210,422,-210</points>
<connection>
<GID>206</GID>
<name>OUT_1</name></connection>
<intersection>422 8</intersection></hsegment></shape></wire>
<wire>
<ID>203 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>448.5,-211.5,456,-211.5</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<connection>
<GID>200</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>204 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>456,-217.5,456,-213.5</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<connection>
<GID>205</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>205 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>448,-223.5,450,-223.5</points>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>449.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>449.5,-223.5,449.5,-218.5</points>
<intersection>-223.5 1</intersection>
<intersection>-218.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>449.5,-218.5,450,-218.5</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>449.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>206 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>449,-221.5,449,-216.5</points>
<intersection>-221.5 23</intersection>
<intersection>-216.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>448.5,-216.5,450,-216.5</points>
<connection>
<GID>196</GID>
<name>OUT</name></connection>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>449 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>449,-221.5,450,-221.5</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>449 0</intersection></hsegment></shape></wire>
<wire>
<ID>207 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>421.5,-196.5,456.5,-196.5</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>421.5 20</intersection>
<intersection>452.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>452.5,-201.5,452.5,-196.5</points>
<intersection>-201.5 16</intersection>
<intersection>-196.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>452.5,-201.5,456.5,-201.5</points>
<connection>
<GID>183</GID>
<name>IN_0</name></connection>
<intersection>452.5 12</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>421.5,-196.5,421.5,-163.5</points>
<intersection>-196.5 1</intersection>
<intersection>-163.5 27</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>404.5,-163.5,421.5,-163.5</points>
<connection>
<GID>207</GID>
<name>OUT_2</name></connection>
<intersection>421.5 20</intersection></hsegment></shape></wire>
<wire>
<ID>208 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>454.5,-198.5,456.5,-198.5</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>454.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>454.5,-203.5,454.5,-198.5</points>
<intersection>-203.5 15</intersection>
<intersection>-198.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>421.5,-203.5,456.5,-203.5</points>
<connection>
<GID>183</GID>
<name>IN_1</name></connection>
<intersection>421.5 17</intersection>
<intersection>454.5 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>421.5,-208,421.5,-203.5</points>
<intersection>-208 18</intersection>
<intersection>-203.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>404.5,-208,421.5,-208</points>
<connection>
<GID>206</GID>
<name>OUT_2</name></connection>
<intersection>421.5 17</intersection></hsegment></shape></wire>
<wire>
<ID>209 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>462.5,-197.5,470,-197.5</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<connection>
<GID>190</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>210 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>470,-203.5,470,-199.5</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<connection>
<GID>189</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>211 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>462,-209.5,464,-209.5</points>
<connection>
<GID>184</GID>
<name>IN_1</name></connection>
<intersection>462 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>462,-212.5,462,-204.5</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<intersection>-209.5 1</intersection>
<intersection>-204.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>462,-204.5,464,-204.5</points>
<connection>
<GID>189</GID>
<name>IN_1</name></connection>
<intersection>462 12</intersection></hsegment></shape></wire>
<wire>
<ID>212 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>463,-207.5,463,-202.5</points>
<intersection>-207.5 23</intersection>
<intersection>-202.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>462.5,-202.5,464,-202.5</points>
<connection>
<GID>183</GID>
<name>OUT</name></connection>
<connection>
<GID>189</GID>
<name>IN_0</name></connection>
<intersection>463 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>463,-207.5,464,-207.5</points>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>463 0</intersection></hsegment></shape></wire>
<wire>
<ID>213 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>468.5,-185.5,471.5,-185.5</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>468.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>468.5,-190.5,468.5,-185.5</points>
<intersection>-190.5 4</intersection>
<intersection>-185.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>420,-190.5,471.5,-190.5</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>420 9</intersection>
<intersection>468.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>420,-190.5,420,-161.5</points>
<intersection>-190.5 4</intersection>
<intersection>-161.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>404.5,-161.5,420,-161.5</points>
<connection>
<GID>207</GID>
<name>OUT_3</name></connection>
<intersection>420 9</intersection></hsegment></shape></wire>
<wire>
<ID>214 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>470,-192.5,470,-187.5</points>
<intersection>-192.5 2</intersection>
<intersection>-187.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>420.5,-192.5,471.5,-192.5</points>
<connection>
<GID>191</GID>
<name>IN_1</name></connection>
<intersection>420.5 8</intersection>
<intersection>470 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>420.5,-206,420.5,-192.5</points>
<intersection>-206 9</intersection>
<intersection>-192.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>404.5,-206,420.5,-206</points>
<connection>
<GID>206</GID>
<name>OUT_3</name></connection>
<intersection>420.5 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>470,-187.5,471.5,-187.5</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<intersection>470 0</intersection></hsegment></shape></wire>
<wire>
<ID>215 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477.5,-186.5,485,-186.5</points>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<connection>
<GID>192</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>216 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>485,-192.5,485,-188.5</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<connection>
<GID>186</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>217 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>476,-198.5,479,-198.5</points>
<connection>
<GID>188</GID>
<name>OUT</name></connection>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<intersection>476 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>476,-198.5,476,-193.5</points>
<intersection>-198.5 1</intersection>
<intersection>-193.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>476,-193.5,479,-193.5</points>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>476 3</intersection></hsegment></shape></wire>
<wire>
<ID>218 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>477.5,-196.5,477.5,-191.5</points>
<connection>
<GID>191</GID>
<name>OUT</name></connection>
<intersection>-196.5 23</intersection>
<intersection>-191.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>477.5,-191.5,479,-191.5</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>477.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>477.5,-196.5,479,-196.5</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>477.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>496.5,-233.5,496.5,-187</points>
<intersection>-233.5 2</intersection>
<intersection>-187 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>496.5,-187,500.5,-187</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>496.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>442,-233.5,496.5,-233.5</points>
<connection>
<GID>204</GID>
<name>OUT</name></connection>
<intersection>496.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>495.5,-222.5,495.5,-186</points>
<intersection>-222.5 2</intersection>
<intersection>-186 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>495.5,-186,500.5,-186</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>495.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>456,-222.5,495.5,-222.5</points>
<connection>
<GID>194</GID>
<name>OUT</name></connection>
<intersection>495.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>221 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>494.5,-208.5,494.5,-185</points>
<intersection>-208.5 2</intersection>
<intersection>-185 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>494.5,-185,500.5,-185</points>
<connection>
<GID>199</GID>
<name>IN_2</name></connection>
<intersection>494.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>470,-208.5,494.5,-208.5</points>
<connection>
<GID>184</GID>
<name>OUT</name></connection>
<intersection>494.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>222 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>493.5,-197.5,493.5,-184</points>
<intersection>-197.5 2</intersection>
<intersection>-184 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>493.5,-184,500.5,-184</points>
<connection>
<GID>199</GID>
<name>IN_3</name></connection>
<intersection>493.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>485,-197.5,493.5,-197.5</points>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<intersection>493.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>223 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>442,-183,500.5,-183</points>
<connection>
<GID>199</GID>
<name>IN_4</name></connection>
<intersection>442 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>442,-183,442,-181.5</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>-183 1</intersection></vsegment></shape></wire>
<wire>
<ID>224 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>493.5,-182,493.5,-170.5</points>
<intersection>-182 1</intersection>
<intersection>-170.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>493.5,-182,500.5,-182</points>
<connection>
<GID>199</GID>
<name>IN_5</name></connection>
<intersection>493.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>456,-170.5,493.5,-170.5</points>
<connection>
<GID>172</GID>
<name>OUT</name></connection>
<intersection>493.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>226 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>495.5,-180,495.5,-145.5</points>
<intersection>-180 1</intersection>
<intersection>-145.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>495.5,-180,500.5,-180</points>
<connection>
<GID>199</GID>
<name>IN_7</name></connection>
<intersection>495.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>485,-145.5,495.5,-145.5</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<intersection>495.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>228 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>423.5,-278.5,428,-278.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>423.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>423.5,-283.5,423.5,-263.5</points>
<intersection>-283.5 16</intersection>
<intersection>-278.5 1</intersection>
<intersection>-263.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>404,-263.5,423.5,-263.5</points>
<connection>
<GID>219</GID>
<name>OUT_0</name></connection>
<intersection>423.5 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>423.5,-283.5,428,-283.5</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>423.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>229 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>422.5,-280.5,428,-280.5</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>422.5 4</intersection>
<intersection>425.5 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>422.5,-308,422.5,-280.5</points>
<intersection>-308 14</intersection>
<intersection>-280.5 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>425.5,-285.5,425.5,-280.5</points>
<intersection>-285.5 15</intersection>
<intersection>-280.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>404,-308,422.5,-308</points>
<connection>
<GID>211</GID>
<name>OUT_0</name></connection>
<intersection>422.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>425.5,-285.5,428,-285.5</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>425.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>230 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>434,-279.5,441.5,-279.5</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<connection>
<GID>214</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>231 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>441.5,-285.5,441.5,-281.5</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<connection>
<GID>216</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>232 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>432,-293,492,-293</points>
<intersection>432 12</intersection>
<intersection>435.5 19</intersection>
<intersection>492 15</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>432,-293,432,-286.5</points>
<intersection>-293 1</intersection>
<intersection>-286.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>432,-286.5,435.5,-286.5</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>432 12</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>492,-296.5,492,-293</points>
<intersection>-296.5 32</intersection>
<intersection>-293 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>435.5,-293,435.5,-291.5</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>-293 1</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>490.5,-296.5,492,-296.5</points>
<connection>
<GID>239</GID>
<name>OUT</name></connection>
<intersection>492 15</intersection></hsegment></shape></wire>
<wire>
<ID>233 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434,-289.5,434,-284.5</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<intersection>-289.5 23</intersection>
<intersection>-284.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>434,-284.5,435.5,-284.5</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>434 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>434,-289.5,435.5,-289.5</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>434 0</intersection></hsegment></shape></wire>
<wire>
<ID>234 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>404,-261.5,442,-261.5</points>
<connection>
<GID>219</GID>
<name>OUT_1</name></connection>
<intersection>442 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>442,-272.5,442,-261.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>-261.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>235 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>440,-274.5,440,-269.5</points>
<intersection>-274.5 2</intersection>
<intersection>-269.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>421.5,-274.5,442,-274.5</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<intersection>421.5 8</intersection>
<intersection>440 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>440,-269.5,442,-269.5</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>440 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>421.5,-306,421.5,-274.5</points>
<intersection>-306 9</intersection>
<intersection>-274.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>404,-306,421.5,-306</points>
<connection>
<GID>211</GID>
<name>OUT_1</name></connection>
<intersection>421.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>236 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>448,-268.5,455.5,-268.5</points>
<connection>
<GID>231</GID>
<name>OUT</name></connection>
<connection>
<GID>218</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>237 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>455.5,-274.5,455.5,-270.5</points>
<connection>
<GID>212</GID>
<name>OUT</name></connection>
<connection>
<GID>218</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>238 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>447.5,-280.5,449.5,-280.5</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<intersection>447.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>447.5,-280.5,447.5,-275.5</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>-280.5 1</intersection>
<intersection>-275.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>447.5,-275.5,449.5,-275.5</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<intersection>447.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>239 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>448,-278.5,448,-273.5</points>
<connection>
<GID>223</GID>
<name>OUT</name></connection>
<intersection>-278.5 23</intersection>
<intersection>-273.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>448,-273.5,449.5,-273.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<intersection>448 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>448,-278.5,449.5,-278.5</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>448 0</intersection></hsegment></shape></wire>
<wire>
<ID>240 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>404,-259.5,456,-259.5</points>
<connection>
<GID>219</GID>
<name>OUT_2</name></connection>
<intersection>451 20</intersection>
<intersection>456 23</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>451,-259.5,451,-253.5</points>
<intersection>-259.5 1</intersection>
<intersection>-253.5 22</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>451,-253.5,456,-253.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>451 20</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>456,-259.5,456,-258.5</points>
<connection>
<GID>235</GID>
<name>IN_0</name></connection>
<intersection>-259.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>241 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>454,-255.5,456,-255.5</points>
<connection>
<GID>228</GID>
<name>IN_1</name></connection>
<intersection>454 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>454,-260.5,454,-255.5</points>
<intersection>-260.5 15</intersection>
<intersection>-255.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>420.5,-260.5,456,-260.5</points>
<connection>
<GID>235</GID>
<name>IN_1</name></connection>
<intersection>420.5 17</intersection>
<intersection>454 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>420.5,-304,420.5,-260.5</points>
<intersection>-304 18</intersection>
<intersection>-260.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>404,-304,420.5,-304</points>
<connection>
<GID>211</GID>
<name>OUT_2</name></connection>
<intersection>420.5 17</intersection></hsegment></shape></wire>
<wire>
<ID>242 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>462,-254.5,469.5,-254.5</points>
<connection>
<GID>228</GID>
<name>OUT</name></connection>
<connection>
<GID>230</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>243 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>469.5,-260.5,469.5,-256.5</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<connection>
<GID>230</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>244 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>461.5,-266.5,463.5,-266.5</points>
<connection>
<GID>234</GID>
<name>IN_1</name></connection>
<intersection>461.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>461.5,-269.5,461.5,-261.5</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<intersection>-266.5 1</intersection>
<intersection>-261.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>461.5,-261.5,463.5,-261.5</points>
<connection>
<GID>229</GID>
<name>IN_1</name></connection>
<intersection>461.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>245 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>462,-264.5,462,-259.5</points>
<connection>
<GID>235</GID>
<name>OUT</name></connection>
<intersection>-264.5 23</intersection>
<intersection>-259.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>462,-259.5,463.5,-259.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>462 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>462,-264.5,463.5,-264.5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<intersection>462 0</intersection></hsegment></shape></wire>
<wire>
<ID>246 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>419.5,-242.5,471,-242.5</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>419.5 6</intersection>
<intersection>468.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>468.5,-247.5,468.5,-242.5</points>
<intersection>-247.5 4</intersection>
<intersection>-242.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>468.5,-247.5,471,-247.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>468.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>419.5,-257.5,419.5,-242.5</points>
<intersection>-257.5 8</intersection>
<intersection>-242.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>404,-257.5,419.5,-257.5</points>
<connection>
<GID>219</GID>
<name>OUT_3</name></connection>
<intersection>419.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>247 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>469.5,-249.5,469.5,-244.5</points>
<intersection>-249.5 2</intersection>
<intersection>-244.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>420,-249.5,471,-249.5</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<intersection>420 8</intersection>
<intersection>469.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>420,-302,420,-249.5</points>
<intersection>-302 9</intersection>
<intersection>-249.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>404,-302,420,-302</points>
<connection>
<GID>211</GID>
<name>OUT_3</name></connection>
<intersection>420 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>469.5,-244.5,471,-244.5</points>
<connection>
<GID>226</GID>
<name>IN_1</name></connection>
<intersection>469.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>248 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>477,-243.5,484.5,-243.5</points>
<connection>
<GID>226</GID>
<name>OUT</name></connection>
<connection>
<GID>232</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>249 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>484.5,-249.5,484.5,-245.5</points>
<connection>
<GID>232</GID>
<name>IN_1</name></connection>
<connection>
<GID>233</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>250 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>475.5,-255.5,478.5,-255.5</points>
<connection>
<GID>230</GID>
<name>OUT</name></connection>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<intersection>477 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>477,-255.5,477,-250.5</points>
<intersection>-255.5 1</intersection>
<intersection>-250.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>477,-250.5,478.5,-250.5</points>
<connection>
<GID>233</GID>
<name>IN_1</name></connection>
<intersection>477 3</intersection></hsegment></shape></wire>
<wire>
<ID>251 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>477,-253.5,477,-248.5</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<intersection>-253.5 23</intersection>
<intersection>-248.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>477,-248.5,478.5,-248.5</points>
<connection>
<GID>233</GID>
<name>IN_0</name></connection>
<intersection>477 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>477,-253.5,478.5,-253.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>477 0</intersection></hsegment></shape></wire>
<wire>
<ID>252 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>423.5,-330.5,428,-330.5</points>
<connection>
<GID>250</GID>
<name>IN_0</name></connection>
<intersection>423.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>423.5,-335.5,423.5,-276.5</points>
<intersection>-335.5 16</intersection>
<intersection>-330.5 1</intersection>
<intersection>-276.5 24</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>423.5,-335.5,428,-335.5</points>
<connection>
<GID>255</GID>
<name>IN_0</name></connection>
<intersection>423.5 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>404,-276.5,423.5,-276.5</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<intersection>423.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>253 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>422.5,-332.5,428,-332.5</points>
<connection>
<GID>250</GID>
<name>IN_1</name></connection>
<intersection>422.5 4</intersection>
<intersection>425.5 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>422.5,-332.5,422.5,-321</points>
<intersection>-332.5 2</intersection>
<intersection>-321 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>425.5,-337.5,425.5,-332.5</points>
<intersection>-337.5 15</intersection>
<intersection>-332.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>404,-321,422.5,-321</points>
<connection>
<GID>259</GID>
<name>OUT_0</name></connection>
<intersection>422.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>425.5,-337.5,428,-337.5</points>
<connection>
<GID>255</GID>
<name>IN_1</name></connection>
<intersection>425.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>254 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>434,-331.5,441.5,-331.5</points>
<connection>
<GID>250</GID>
<name>OUT</name></connection>
<connection>
<GID>256</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>255 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>441.5,-337.5,441.5,-333.5</points>
<connection>
<GID>254</GID>
<name>OUT</name></connection>
<connection>
<GID>256</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>256 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>404,-343.5,435.5,-343.5</points>
<connection>
<GID>251</GID>
<name>OUT_0</name></connection>
<connection>
<GID>257</GID>
<name>IN_1</name></connection>
<intersection>433 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>433,-343.5,433,-338.5</points>
<intersection>-343.5 1</intersection>
<intersection>-338.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>433,-338.5,435.5,-338.5</points>
<connection>
<GID>254</GID>
<name>IN_1</name></connection>
<intersection>433 12</intersection></hsegment></shape></wire>
<wire>
<ID>257 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>434,-341.5,434,-336.5</points>
<connection>
<GID>255</GID>
<name>OUT</name></connection>
<intersection>-341.5 23</intersection>
<intersection>-336.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>434,-336.5,435.5,-336.5</points>
<connection>
<GID>254</GID>
<name>IN_0</name></connection>
<intersection>434 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>434,-341.5,435.5,-341.5</points>
<connection>
<GID>257</GID>
<name>IN_0</name></connection>
<intersection>434 0</intersection></hsegment></shape></wire>
<wire>
<ID>315 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>545.5,-210.5,565.5,-210.5</points>
<connection>
<GID>331</GID>
<name>IN_0</name></connection>
<intersection>545.5 6</intersection>
<intersection>562.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>562.5,-215.5,562.5,-210.5</points>
<intersection>-215.5 4</intersection>
<intersection>-210.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>562.5,-215.5,565.5,-215.5</points>
<connection>
<GID>323</GID>
<name>IN_0</name></connection>
<intersection>562.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>545.5,-210.5,545.5,-165.5</points>
<intersection>-210.5 1</intersection>
<intersection>-165.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>527.5,-165.5,545.5,-165.5</points>
<connection>
<GID>313</GID>
<name>OUT_1</name></connection>
<intersection>545.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>316 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>563.5,-217.5,563.5,-212.5</points>
<intersection>-217.5 2</intersection>
<intersection>-212.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>545,-217.5,565.5,-217.5</points>
<connection>
<GID>323</GID>
<name>IN_1</name></connection>
<intersection>545 8</intersection>
<intersection>563.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>563.5,-212.5,565.5,-212.5</points>
<connection>
<GID>331</GID>
<name>IN_1</name></connection>
<intersection>563.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>545,-217.5,545,-210</points>
<intersection>-217.5 2</intersection>
<intersection>-210 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>527.5,-210,545,-210</points>
<connection>
<GID>314</GID>
<name>OUT_1</name></connection>
<intersection>545 8</intersection></hsegment></shape></wire>
<wire>
<ID>317 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>571.5,-211.5,579,-211.5</points>
<connection>
<GID>331</GID>
<name>OUT</name></connection>
<connection>
<GID>320</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>318 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>579,-217.5,579,-213.5</points>
<connection>
<GID>320</GID>
<name>IN_1</name></connection>
<connection>
<GID>315</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>319 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>571,-223.5,573,-223.5</points>
<connection>
<GID>325</GID>
<name>IN_1</name></connection>
<connection>
<GID>317</GID>
<name>OUT</name></connection>
<intersection>572.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>572.5,-223.5,572.5,-218.5</points>
<intersection>-223.5 1</intersection>
<intersection>-218.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>572.5,-218.5,573,-218.5</points>
<connection>
<GID>315</GID>
<name>IN_1</name></connection>
<intersection>572.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>320 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>572,-221.5,572,-216.5</points>
<intersection>-221.5 23</intersection>
<intersection>-216.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>571.5,-216.5,573,-216.5</points>
<connection>
<GID>323</GID>
<name>OUT</name></connection>
<connection>
<GID>315</GID>
<name>IN_0</name></connection>
<intersection>572 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>572,-221.5,573,-221.5</points>
<connection>
<GID>325</GID>
<name>IN_0</name></connection>
<intersection>572 0</intersection></hsegment></shape></wire>
<wire>
<ID>321 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>544.5,-196.5,579.5,-196.5</points>
<connection>
<GID>328</GID>
<name>IN_0</name></connection>
<intersection>544.5 20</intersection>
<intersection>575.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>575.5,-201.5,575.5,-196.5</points>
<intersection>-201.5 16</intersection>
<intersection>-196.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>575.5,-201.5,579.5,-201.5</points>
<connection>
<GID>335</GID>
<name>IN_0</name></connection>
<intersection>575.5 12</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>544.5,-196.5,544.5,-163.5</points>
<intersection>-196.5 1</intersection>
<intersection>-163.5 27</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>527.5,-163.5,544.5,-163.5</points>
<connection>
<GID>313</GID>
<name>OUT_2</name></connection>
<intersection>544.5 20</intersection></hsegment></shape></wire>
<wire>
<ID>322 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>577.5,-198.5,579.5,-198.5</points>
<connection>
<GID>328</GID>
<name>IN_1</name></connection>
<intersection>577.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>577.5,-203.5,577.5,-198.5</points>
<intersection>-203.5 15</intersection>
<intersection>-198.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>544.5,-203.5,579.5,-203.5</points>
<connection>
<GID>335</GID>
<name>IN_1</name></connection>
<intersection>544.5 17</intersection>
<intersection>577.5 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>544.5,-208,544.5,-203.5</points>
<intersection>-208 18</intersection>
<intersection>-203.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>527.5,-208,544.5,-208</points>
<connection>
<GID>314</GID>
<name>OUT_2</name></connection>
<intersection>544.5 17</intersection></hsegment></shape></wire>
<wire>
<ID>323 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585.5,-197.5,593,-197.5</points>
<connection>
<GID>330</GID>
<name>IN_0</name></connection>
<connection>
<GID>328</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>324 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>593,-203.5,593,-199.5</points>
<connection>
<GID>330</GID>
<name>IN_1</name></connection>
<connection>
<GID>329</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>325 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-209.5,587,-209.5</points>
<connection>
<GID>334</GID>
<name>IN_1</name></connection>
<intersection>585 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>585,-212.5,585,-204.5</points>
<connection>
<GID>320</GID>
<name>OUT</name></connection>
<intersection>-209.5 1</intersection>
<intersection>-204.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>585,-204.5,587,-204.5</points>
<connection>
<GID>329</GID>
<name>IN_1</name></connection>
<intersection>585 12</intersection></hsegment></shape></wire>
<wire>
<ID>326 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>586,-207.5,586,-202.5</points>
<intersection>-207.5 23</intersection>
<intersection>-202.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>585.5,-202.5,587,-202.5</points>
<connection>
<GID>335</GID>
<name>OUT</name></connection>
<connection>
<GID>329</GID>
<name>IN_0</name></connection>
<intersection>586 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>586,-207.5,587,-207.5</points>
<connection>
<GID>334</GID>
<name>IN_0</name></connection>
<intersection>586 0</intersection></hsegment></shape></wire>
<wire>
<ID>327 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>591.5,-185.5,594.5,-185.5</points>
<connection>
<GID>326</GID>
<name>IN_0</name></connection>
<intersection>591.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>591.5,-190.5,591.5,-185.5</points>
<intersection>-190.5 4</intersection>
<intersection>-185.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>543,-190.5,594.5,-190.5</points>
<connection>
<GID>327</GID>
<name>IN_0</name></connection>
<intersection>543 9</intersection>
<intersection>591.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>543,-190.5,543,-161.5</points>
<intersection>-190.5 4</intersection>
<intersection>-161.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>527.5,-161.5,543,-161.5</points>
<connection>
<GID>313</GID>
<name>OUT_3</name></connection>
<intersection>543 9</intersection></hsegment></shape></wire>
<wire>
<ID>328 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>593,-192.5,593,-187.5</points>
<intersection>-192.5 2</intersection>
<intersection>-187.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>543.5,-192.5,594.5,-192.5</points>
<connection>
<GID>327</GID>
<name>IN_1</name></connection>
<intersection>543.5 8</intersection>
<intersection>593 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>543.5,-206,543.5,-192.5</points>
<intersection>-206 9</intersection>
<intersection>-192.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>527.5,-206,543.5,-206</points>
<connection>
<GID>314</GID>
<name>OUT_3</name></connection>
<intersection>543.5 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>593,-187.5,594.5,-187.5</points>
<connection>
<GID>326</GID>
<name>IN_1</name></connection>
<intersection>593 0</intersection></hsegment></shape></wire>
<wire>
<ID>329 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600.5,-186.5,608,-186.5</points>
<connection>
<GID>332</GID>
<name>IN_0</name></connection>
<connection>
<GID>326</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>330 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>608,-192.5,608,-188.5</points>
<connection>
<GID>333</GID>
<name>OUT</name></connection>
<connection>
<GID>332</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>331 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>599,-198.5,602,-198.5</points>
<connection>
<GID>324</GID>
<name>IN_1</name></connection>
<intersection>599 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>599,-198.5,599,-193.5</points>
<connection>
<GID>330</GID>
<name>OUT</name></connection>
<intersection>-198.5 1</intersection>
<intersection>-193.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>599,-193.5,602,-193.5</points>
<connection>
<GID>333</GID>
<name>IN_1</name></connection>
<intersection>599 3</intersection></hsegment></shape></wire>
<wire>
<ID>332 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>600.5,-196.5,600.5,-191.5</points>
<connection>
<GID>327</GID>
<name>OUT</name></connection>
<intersection>-196.5 23</intersection>
<intersection>-191.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>600.5,-191.5,602,-191.5</points>
<connection>
<GID>333</GID>
<name>IN_0</name></connection>
<intersection>600.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>600.5,-196.5,602,-196.5</points>
<connection>
<GID>324</GID>
<name>IN_0</name></connection>
<intersection>600.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>333 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>619.5,-233.5,619.5,-186.5</points>
<intersection>-233.5 2</intersection>
<intersection>-186.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>619.5,-186.5,642,-186.5</points>
<connection>
<GID>321</GID>
<name>IN_0</name></connection>
<intersection>619.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>565,-233.5,619.5,-233.5</points>
<connection>
<GID>316</GID>
<name>OUT</name></connection>
<intersection>619.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>334 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,-222.5,618.5,-185.5</points>
<intersection>-222.5 2</intersection>
<intersection>-185.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618.5,-185.5,642,-185.5</points>
<connection>
<GID>321</GID>
<name>IN_1</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>579,-222.5,618.5,-222.5</points>
<connection>
<GID>325</GID>
<name>OUT</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>335 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>617.5,-208.5,617.5,-184.5</points>
<intersection>-208.5 2</intersection>
<intersection>-184.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>617.5,-184.5,642,-184.5</points>
<connection>
<GID>321</GID>
<name>IN_2</name></connection>
<intersection>617.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>593,-208.5,617.5,-208.5</points>
<connection>
<GID>334</GID>
<name>OUT</name></connection>
<intersection>617.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>336 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>616.5,-197.5,616.5,-183.5</points>
<intersection>-197.5 2</intersection>
<intersection>-183.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,-183.5,642,-183.5</points>
<connection>
<GID>321</GID>
<name>IN_3</name></connection>
<intersection>616.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>608,-197.5,616.5,-197.5</points>
<connection>
<GID>324</GID>
<name>OUT</name></connection>
<intersection>616.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>337 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>565,-182.5,642,-182.5</points>
<connection>
<GID>321</GID>
<name>IN_4</name></connection>
<intersection>565 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>565,-182.5,565,-181.5</points>
<connection>
<GID>358</GID>
<name>OUT</name></connection>
<intersection>-182.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>338 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>616.5,-181.5,616.5,-170.5</points>
<intersection>-181.5 1</intersection>
<intersection>-170.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>616.5,-181.5,642,-181.5</points>
<connection>
<GID>321</GID>
<name>IN_5</name></connection>
<intersection>616.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>579,-170.5,616.5,-170.5</points>
<connection>
<GID>346</GID>
<name>OUT</name></connection>
<intersection>616.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>339 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>617.5,-180.5,617.5,-156.5</points>
<intersection>-180.5 1</intersection>
<intersection>-156.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>617.5,-180.5,642,-180.5</points>
<connection>
<GID>321</GID>
<name>IN_6</name></connection>
<intersection>617.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>593,-156.5,617.5,-156.5</points>
<connection>
<GID>337</GID>
<name>OUT</name></connection>
<intersection>617.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>340 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>618.5,-179.5,618.5,-145.5</points>
<intersection>-179.5 1</intersection>
<intersection>-145.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>618.5,-179.5,642,-179.5</points>
<connection>
<GID>321</GID>
<name>IN_7</name></connection>
<intersection>618.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>608,-145.5,618.5,-145.5</points>
<connection>
<GID>347</GID>
<name>OUT</name></connection>
<intersection>618.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>341 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>619.5,-177,619.5,-135.5</points>
<intersection>-177 1</intersection>
<intersection>-135.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>619.5,-177,642,-177</points>
<connection>
<GID>312</GID>
<name>IN_0</name></connection>
<intersection>619.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>614,-135.5,619.5,-135.5</points>
<connection>
<GID>339</GID>
<name>OUT</name></connection>
<intersection>619.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>342 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>546.5,-278.5,551,-278.5</points>
<connection>
<GID>300</GID>
<name>IN_0</name></connection>
<intersection>546.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>546.5,-283.5,546.5,-263.5</points>
<intersection>-283.5 16</intersection>
<intersection>-278.5 1</intersection>
<intersection>-263.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>527,-263.5,546.5,-263.5</points>
<connection>
<GID>301</GID>
<name>OUT_0</name></connection>
<intersection>546.5 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>546.5,-283.5,551,-283.5</points>
<connection>
<GID>305</GID>
<name>IN_0</name></connection>
<intersection>546.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>343 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>545.5,-280.5,551,-280.5</points>
<connection>
<GID>300</GID>
<name>IN_1</name></connection>
<intersection>545.5 4</intersection>
<intersection>548.5 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>545.5,-308,545.5,-280.5</points>
<intersection>-308 14</intersection>
<intersection>-280.5 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>548.5,-285.5,548.5,-280.5</points>
<intersection>-285.5 15</intersection>
<intersection>-280.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>527,-308,545.5,-308</points>
<connection>
<GID>309</GID>
<name>OUT_0</name></connection>
<intersection>545.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>548.5,-285.5,551,-285.5</points>
<connection>
<GID>305</GID>
<name>IN_1</name></connection>
<intersection>548.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>344 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>557,-279.5,564.5,-279.5</points>
<connection>
<GID>300</GID>
<name>OUT</name></connection>
<connection>
<GID>306</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>345 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>564.5,-285.5,564.5,-281.5</points>
<connection>
<GID>304</GID>
<name>OUT</name></connection>
<connection>
<GID>306</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>346 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>555,-293,615,-293</points>
<intersection>555 12</intersection>
<intersection>558.5 19</intersection>
<intersection>615 15</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>555,-293,555,-286.5</points>
<intersection>-293 1</intersection>
<intersection>-286.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>555,-286.5,558.5,-286.5</points>
<connection>
<GID>304</GID>
<name>IN_1</name></connection>
<intersection>555 12</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>615,-296.5,615,-293</points>
<intersection>-296.5 32</intersection>
<intersection>-293 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>558.5,-293,558.5,-291.5</points>
<connection>
<GID>307</GID>
<name>IN_1</name></connection>
<intersection>-293 1</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>613.5,-296.5,615,-296.5</points>
<connection>
<GID>282</GID>
<name>OUT</name></connection>
<intersection>615 15</intersection></hsegment></shape></wire>
<wire>
<ID>347 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>557,-289.5,557,-284.5</points>
<connection>
<GID>305</GID>
<name>OUT</name></connection>
<intersection>-289.5 23</intersection>
<intersection>-284.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>557,-284.5,558.5,-284.5</points>
<connection>
<GID>304</GID>
<name>IN_0</name></connection>
<intersection>557 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>557,-289.5,558.5,-289.5</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>557 0</intersection></hsegment></shape></wire>
<wire>
<ID>348 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>527,-261.5,565,-261.5</points>
<connection>
<GID>301</GID>
<name>OUT_1</name></connection>
<intersection>565 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>565,-272.5,565,-261.5</points>
<connection>
<GID>290</GID>
<name>IN_0</name></connection>
<connection>
<GID>298</GID>
<name>IN_0</name></connection>
<intersection>-261.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>349 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>563,-274.5,563,-269.5</points>
<intersection>-274.5 2</intersection>
<intersection>-269.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>544.5,-274.5,565,-274.5</points>
<connection>
<GID>298</GID>
<name>IN_1</name></connection>
<intersection>544.5 8</intersection>
<intersection>563 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>563,-269.5,565,-269.5</points>
<connection>
<GID>290</GID>
<name>IN_1</name></connection>
<intersection>563 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>544.5,-306,544.5,-274.5</points>
<intersection>-306 9</intersection>
<intersection>-274.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>527,-306,544.5,-306</points>
<connection>
<GID>309</GID>
<name>OUT_1</name></connection>
<intersection>544.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>350 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>571,-268.5,578.5,-268.5</points>
<connection>
<GID>290</GID>
<name>OUT</name></connection>
<connection>
<GID>302</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>351 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>578.5,-274.5,578.5,-270.5</points>
<connection>
<GID>302</GID>
<name>IN_1</name></connection>
<connection>
<GID>308</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>352 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>570.5,-280.5,572.5,-280.5</points>
<connection>
<GID>296</GID>
<name>IN_1</name></connection>
<intersection>570.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>570.5,-280.5,570.5,-275.5</points>
<connection>
<GID>306</GID>
<name>OUT</name></connection>
<intersection>-280.5 1</intersection>
<intersection>-275.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>570.5,-275.5,572.5,-275.5</points>
<connection>
<GID>308</GID>
<name>IN_1</name></connection>
<intersection>570.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>353 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>571,-278.5,571,-273.5</points>
<connection>
<GID>298</GID>
<name>OUT</name></connection>
<intersection>-278.5 23</intersection>
<intersection>-273.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>571,-273.5,572.5,-273.5</points>
<connection>
<GID>308</GID>
<name>IN_0</name></connection>
<intersection>571 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>571,-278.5,572.5,-278.5</points>
<connection>
<GID>296</GID>
<name>IN_0</name></connection>
<intersection>571 0</intersection></hsegment></shape></wire>
<wire>
<ID>354 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>527,-259.5,579,-259.5</points>
<connection>
<GID>301</GID>
<name>OUT_2</name></connection>
<intersection>574 20</intersection>
<intersection>579 23</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>574,-259.5,574,-253.5</points>
<intersection>-259.5 1</intersection>
<intersection>-253.5 22</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>574,-253.5,579,-253.5</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>574 20</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>579,-259.5,579,-258.5</points>
<connection>
<GID>286</GID>
<name>IN_0</name></connection>
<intersection>-259.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>355 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>577,-255.5,579,-255.5</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<intersection>577 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>577,-260.5,577,-255.5</points>
<intersection>-260.5 15</intersection>
<intersection>-255.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>543.5,-260.5,579,-260.5</points>
<connection>
<GID>286</GID>
<name>IN_1</name></connection>
<intersection>543.5 17</intersection>
<intersection>577 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>543.5,-304,543.5,-260.5</points>
<intersection>-304 18</intersection>
<intersection>-260.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>527,-304,543.5,-304</points>
<connection>
<GID>309</GID>
<name>OUT_2</name></connection>
<intersection>543.5 17</intersection></hsegment></shape></wire>
<wire>
<ID>356 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>585,-254.5,592.5,-254.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<connection>
<GID>293</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>357 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-260.5,592.5,-256.5</points>
<connection>
<GID>291</GID>
<name>IN_1</name></connection>
<connection>
<GID>292</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>358 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>584.5,-266.5,586.5,-266.5</points>
<connection>
<GID>287</GID>
<name>IN_1</name></connection>
<intersection>584.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>584.5,-269.5,584.5,-261.5</points>
<connection>
<GID>302</GID>
<name>OUT</name></connection>
<intersection>-266.5 1</intersection>
<intersection>-261.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>584.5,-261.5,586.5,-261.5</points>
<connection>
<GID>292</GID>
<name>IN_1</name></connection>
<intersection>584.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>359 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>585,-264.5,585,-259.5</points>
<connection>
<GID>286</GID>
<name>OUT</name></connection>
<intersection>-264.5 23</intersection>
<intersection>-259.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>585,-259.5,586.5,-259.5</points>
<connection>
<GID>292</GID>
<name>IN_0</name></connection>
<intersection>585 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>585,-264.5,586.5,-264.5</points>
<connection>
<GID>287</GID>
<name>IN_0</name></connection>
<intersection>585 0</intersection></hsegment></shape></wire>
<wire>
<ID>360 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>542.5,-242.5,594,-242.5</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>542.5 6</intersection>
<intersection>591.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>591.5,-247.5,591.5,-242.5</points>
<intersection>-247.5 4</intersection>
<intersection>-242.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>591.5,-247.5,594,-247.5</points>
<connection>
<GID>294</GID>
<name>IN_0</name></connection>
<intersection>591.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>542.5,-257.5,542.5,-242.5</points>
<intersection>-257.5 8</intersection>
<intersection>-242.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>527,-257.5,542.5,-257.5</points>
<connection>
<GID>301</GID>
<name>OUT_3</name></connection>
<intersection>542.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>361 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>592.5,-249.5,592.5,-244.5</points>
<intersection>-249.5 2</intersection>
<intersection>-244.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>543,-249.5,594,-249.5</points>
<connection>
<GID>294</GID>
<name>IN_1</name></connection>
<intersection>543 8</intersection>
<intersection>592.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>543,-302,543,-249.5</points>
<intersection>-302 9</intersection>
<intersection>-249.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>527,-302,543,-302</points>
<connection>
<GID>309</GID>
<name>OUT_3</name></connection>
<intersection>543 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>592.5,-244.5,594,-244.5</points>
<connection>
<GID>295</GID>
<name>IN_1</name></connection>
<intersection>592.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>362 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>600,-243.5,607.5,-243.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<connection>
<GID>295</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>363 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>607.5,-249.5,607.5,-245.5</points>
<connection>
<GID>288</GID>
<name>OUT</name></connection>
<connection>
<GID>289</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>364 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>598.5,-255.5,601.5,-255.5</points>
<connection>
<GID>291</GID>
<name>OUT</name></connection>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>599 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>599,-255.5,599,-250.5</points>
<intersection>-255.5 1</intersection>
<intersection>-250.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>599,-250.5,601.5,-250.5</points>
<connection>
<GID>288</GID>
<name>IN_1</name></connection>
<intersection>599 3</intersection></hsegment></shape></wire>
<wire>
<ID>365 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>600,-253.5,600,-248.5</points>
<connection>
<GID>294</GID>
<name>OUT</name></connection>
<intersection>-253.5 23</intersection>
<intersection>-248.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>600,-248.5,601.5,-248.5</points>
<connection>
<GID>288</GID>
<name>IN_0</name></connection>
<intersection>600 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>600,-253.5,601.5,-253.5</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>600 0</intersection></hsegment></shape></wire>
<wire>
<ID>366 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>546.5,-330.5,551,-330.5</points>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>546.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>546.5,-335.5,546.5,-276.5</points>
<intersection>-335.5 16</intersection>
<intersection>-330.5 1</intersection>
<intersection>-276.5 24</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>546.5,-335.5,551,-335.5</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>546.5 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>527,-276.5,546.5,-276.5</points>
<connection>
<GID>363</GID>
<name>OUT_0</name></connection>
<intersection>546.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>367 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>545.5,-332.5,551,-332.5</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<intersection>545.5 4</intersection>
<intersection>548.5 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>545.5,-332.5,545.5,-321</points>
<intersection>-332.5 2</intersection>
<intersection>-321 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>548.5,-337.5,548.5,-332.5</points>
<intersection>-337.5 15</intersection>
<intersection>-332.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>527,-321,545.5,-321</points>
<connection>
<GID>362</GID>
<name>OUT_0</name></connection>
<intersection>545.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>548.5,-337.5,551,-337.5</points>
<connection>
<GID>266</GID>
<name>IN_1</name></connection>
<intersection>548.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>368 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>557,-331.5,564.5,-331.5</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<connection>
<GID>271</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>369 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>564.5,-337.5,564.5,-333.5</points>
<connection>
<GID>265</GID>
<name>IN_1</name></connection>
<connection>
<GID>267</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>370 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>510.5,-343.5,558.5,-343.5</points>
<connection>
<GID>264</GID>
<name>IN_1</name></connection>
<intersection>510.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>510.5,-343.5,510.5,-135.5</points>
<intersection>-343.5 1</intersection>
<intersection>-338.5 14</intersection>
<intersection>-135.5 15</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>510.5,-338.5,558.5,-338.5</points>
<connection>
<GID>267</GID>
<name>IN_1</name></connection>
<intersection>510.5 12</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>491,-135.5,510.5,-135.5</points>
<connection>
<GID>179</GID>
<name>OUT</name></connection>
<intersection>510.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>371 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>557,-341.5,557,-336.5</points>
<connection>
<GID>266</GID>
<name>OUT</name></connection>
<intersection>-341.5 23</intersection>
<intersection>-336.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>557,-336.5,558.5,-336.5</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>557 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>557,-341.5,558.5,-341.5</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>557 0</intersection></hsegment></shape></wire></page 0></circuit>