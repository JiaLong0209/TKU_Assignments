
<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-32.95,39.6893,61.95,-63.2229</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>14.5,-13</position>
<gparam>LABEL_TEXT Go to https://cedar.to/vjyQw7 to download the latest version!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>14.5,-9.5</position>
<gparam>LABEL_TEXT Error: This file was made with a newer version of Cedar Logic!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 0>
</circuit>
<throw_away></throw_away>

	<version>2.3.8 | 2024-10-27 09:03:56</version><circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>96.2489,-109.213,404.698,-273.282</PageViewport>
<gate>
<ID>231</ID>
<type>DD_KEYPAD_HEX</type>
<position>223.5,-222.5</position>
<output>
<ID>OUT_0</ID>172 </output>
<output>
<ID>OUT_1</ID>178 </output>
<output>
<ID>OUT_2</ID>184 </output>
<output>
<ID>OUT_3</ID>190 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>230</ID>
<type>AA_AND2</type>
<position>277,-192</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>180 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>229</ID>
<type>AI_XOR2</type>
<position>263,-208</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>175 </input>
<output>
<ID>OUT</ID>223 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>228</ID>
<type>AE_OR2</type>
<position>269,-198</position>
<input>
<ID>IN_0</ID>173 </input>
<input>
<ID>IN_1</ID>174 </input>
<output>
<ID>OUT</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>AI_XOR2</type>
<position>255.5,-202</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT</ID>176 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>226</ID>
<type>AA_AND2</type>
<position>263,-203</position>
<input>
<ID>IN_0</ID>176 </input>
<input>
<ID>IN_1</ID>175 </input>
<output>
<ID>OUT</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>225</ID>
<type>AA_LABEL</type>
<position>215.5,-235.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>224</ID>
<type>AE_OR2</type>
<position>283,-187</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>180 </input>
<output>
<ID>OUT</ID>187 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>223</ID>
<type>DD_KEYPAD_HEX</type>
<position>223.5,-178</position>
<output>
<ID>OUT_0</ID>171 </output>
<output>
<ID>OUT_1</ID>177 </output>
<output>
<ID>OUT_2</ID>183 </output>
<output>
<ID>OUT_3</ID>189 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_LABEL</type>
<position>274,-156</position>
<gparam>LABEL_TEXT 8-Bits Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>255.5,-197</position>
<input>
<ID>IN_0</ID>171 </input>
<input>
<ID>IN_1</ID>172 </input>
<output>
<ID>OUT</ID>173 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_LABEL</type>
<position>215.5,-178</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AI_XOR2</type>
<position>269.5,-191</position>
<input>
<ID>IN_0</ID>177 </input>
<input>
<ID>IN_1</ID>178 </input>
<output>
<ID>OUT</ID>182 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>218</ID>
<type>AI_XOR2</type>
<position>306,-172</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>193 </input>
<output>
<ID>OUT</ID>226 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>217</ID>
<type>AI_XOR2</type>
<position>277,-197</position>
<input>
<ID>IN_0</ID>182 </input>
<input>
<ID>IN_1</ID>181 </input>
<output>
<ID>OUT</ID>224 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_AND2</type>
<position>298.5,-161</position>
<input>
<ID>IN_0</ID>189 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>191 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>215</ID>
<type>AI_XOR2</type>
<position>298.5,-166</position>
<input>
<ID>IN_0</ID>189 </input>
<input>
<ID>IN_1</ID>190 </input>
<output>
<ID>OUT</ID>194 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_AND2</type>
<position>283.5,-172</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>184 </input>
<output>
<ID>OUT</ID>185 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>213</ID>
<type>AA_AND2</type>
<position>291,-178</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>186 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>212</ID>
<type>AE_OR2</type>
<position>297,-173</position>
<input>
<ID>IN_0</ID>185 </input>
<input>
<ID>IN_1</ID>186 </input>
<output>
<ID>OUT</ID>193 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>211</ID>
<type>AA_AND2</type>
<position>269.5,-186</position>
<input>
<ID>IN_0</ID>177 </input>
<input>
<ID>IN_1</ID>178 </input>
<output>
<ID>OUT</ID>179 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>210</ID>
<type>AE_OR2</type>
<position>312,-162</position>
<input>
<ID>IN_0</ID>191 </input>
<input>
<ID>IN_1</ID>192 </input>
<output>
<ID>OUT</ID>227 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>209</ID>
<type>AA_AND2</type>
<position>306,-167</position>
<input>
<ID>IN_0</ID>194 </input>
<input>
<ID>IN_1</ID>193 </input>
<output>
<ID>OUT</ID>192 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>208</ID>
<type>AI_XOR2</type>
<position>291,-183</position>
<input>
<ID>IN_0</ID>188 </input>
<input>
<ID>IN_1</ID>187 </input>
<output>
<ID>OUT</ID>225 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>AI_XOR2</type>
<position>283.5,-177</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>184 </input>
<output>
<ID>OUT</ID>188 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>206</ID>
<type>AI_XOR2</type>
<position>283.5,-229</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>212 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>AI_XOR2</type>
<position>291,-235</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>221 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>204</ID>
<type>AA_AND2</type>
<position>306,-219</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>216 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>203</ID>
<type>AE_OR2</type>
<position>312,-214</position>
<input>
<ID>IN_0</ID>215 </input>
<input>
<ID>IN_1</ID>216 </input>
<output>
<ID>OUT</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>202</ID>
<type>AA_AND2</type>
<position>269.5,-238</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>202 </input>
<output>
<ID>OUT</ID>203 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>AE_OR2</type>
<position>297,-225</position>
<input>
<ID>IN_0</ID>209 </input>
<input>
<ID>IN_1</ID>210 </input>
<output>
<ID>OUT</ID>217 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>200</ID>
<type>AA_AND2</type>
<position>291,-230</position>
<input>
<ID>IN_0</ID>212 </input>
<input>
<ID>IN_1</ID>211 </input>
<output>
<ID>OUT</ID>210 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>199</ID>
<type>AA_AND2</type>
<position>283.5,-224</position>
<input>
<ID>IN_0</ID>207 </input>
<input>
<ID>IN_1</ID>208 </input>
<output>
<ID>OUT</ID>209 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>198</ID>
<type>AI_XOR2</type>
<position>298.5,-218</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>218 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>197</ID>
<type>AA_AND2</type>
<position>298.5,-213</position>
<input>
<ID>IN_0</ID>213 </input>
<input>
<ID>IN_1</ID>214 </input>
<output>
<ID>OUT</ID>215 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>196</ID>
<type>AA_LABEL</type>
<position>216,-257.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>AI_XOR2</type>
<position>277,-249</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>205 </input>
<output>
<ID>OUT</ID>220 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>194</ID>
<type>AI_XOR2</type>
<position>306,-224</position>
<input>
<ID>IN_0</ID>218 </input>
<input>
<ID>IN_1</ID>217 </input>
<output>
<ID>OUT</ID>222 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>193</ID>
<type>AI_XOR2</type>
<position>269.5,-243</position>
<input>
<ID>IN_0</ID>201 </input>
<input>
<ID>IN_1</ID>202 </input>
<output>
<ID>OUT</ID>206 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>192</ID>
<type>AA_AND2</type>
<position>255.5,-249</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>196 </input>
<output>
<ID>OUT</ID>197 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>191</ID>
<type>DD_KEYPAD_HEX</type>
<position>223.5,-258</position>
<output>
<ID>OUT_0</ID>199 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>190</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>348,-210</position>
<input>
<ID>IN_0</ID>219 </input>
<input>
<ID>IN_1</ID>220 </input>
<input>
<ID>IN_2</ID>221 </input>
<input>
<ID>IN_3</ID>222 </input>
<input>
<ID>IN_4</ID>223 </input>
<input>
<ID>IN_5</ID>224 </input>
<input>
<ID>IN_6</ID>225 </input>
<input>
<ID>IN_7</ID>226 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>189</ID>
<type>AE_OR2</type>
<position>283,-239</position>
<input>
<ID>IN_0</ID>203 </input>
<input>
<ID>IN_1</ID>204 </input>
<output>
<ID>OUT</ID>211 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_AND2</type>
<position>263,-255</position>
<input>
<ID>IN_0</ID>200 </input>
<input>
<ID>IN_1</ID>199 </input>
<output>
<ID>OUT</ID>198 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>187</ID>
<type>AI_XOR2</type>
<position>255.5,-254</position>
<input>
<ID>IN_0</ID>195 </input>
<input>
<ID>IN_1</ID>196 </input>
<output>
<ID>OUT</ID>200 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>186</ID>
<type>AE_OR2</type>
<position>269,-250</position>
<input>
<ID>IN_0</ID>197 </input>
<input>
<ID>IN_1</ID>198 </input>
<output>
<ID>OUT</ID>205 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>185</ID>
<type>AI_XOR2</type>
<position>263,-260</position>
<input>
<ID>IN_0</ID>200 </input>
<input>
<ID>IN_1</ID>199 </input>
<output>
<ID>OUT</ID>219 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>184</ID>
<type>AA_AND2</type>
<position>277,-244</position>
<input>
<ID>IN_0</ID>206 </input>
<input>
<ID>IN_1</ID>205 </input>
<output>
<ID>OUT</ID>204 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>183</ID>
<type>DD_KEYPAD_HEX</type>
<position>223.5,-235.5</position>
<output>
<ID>OUT_0</ID>196 </output>
<output>
<ID>OUT_1</ID>202 </output>
<output>
<ID>OUT_2</ID>208 </output>
<output>
<ID>OUT_3</ID>214 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>182</ID>
<type>DD_KEYPAD_HEX</type>
<position>223.5,-191</position>
<output>
<ID>OUT_0</ID>195 </output>
<output>
<ID>OUT_1</ID>201 </output>
<output>
<ID>OUT_2</ID>207 </output>
<output>
<ID>OUT_3</ID>213 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>181</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>348,-200.5</position>
<input>
<ID>IN_0</ID>227 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>180</ID>
<type>AA_LABEL</type>
<position>215.5,-222.5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>179</ID>
<type>AA_LABEL</type>
<position>215.5,-191.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>AA_LABEL</type>
<position>-71,-204</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>AA_LABEL</type>
<position>-71,-235</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>176</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>61.5,-213</position>
<input>
<ID>IN_0</ID>170 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>175</ID>
<type>DD_KEYPAD_HEX</type>
<position>-63,-203.5</position>
<output>
<ID>OUT_0</ID>138 </output>
<output>
<ID>OUT_1</ID>144 </output>
<output>
<ID>OUT_2</ID>150 </output>
<output>
<ID>OUT_3</ID>156 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>174</ID>
<type>DD_KEYPAD_HEX</type>
<position>-63,-248</position>
<output>
<ID>OUT_0</ID>139 </output>
<output>
<ID>OUT_1</ID>145 </output>
<output>
<ID>OUT_2</ID>151 </output>
<output>
<ID>OUT_3</ID>157 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>173</ID>
<type>AA_AND2</type>
<position>-9.5,-256.5</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>172</ID>
<type>AI_XOR2</type>
<position>-23.5,-272.5</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>162 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>171</ID>
<type>AE_OR2</type>
<position>-17.5,-262.5</position>
<input>
<ID>IN_0</ID>140 </input>
<input>
<ID>IN_1</ID>141 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>170</ID>
<type>AI_XOR2</type>
<position>-31,-266.5</position>
<input>
<ID>IN_0</ID>138 </input>
<input>
<ID>IN_1</ID>139 </input>
<output>
<ID>OUT</ID>143 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>AA_AND2</type>
<position>-23.5,-267.5</position>
<input>
<ID>IN_0</ID>143 </input>
<input>
<ID>IN_1</ID>142 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>167</ID>
<type>AE_OR2</type>
<position>-3.5,-251.5</position>
<input>
<ID>IN_0</ID>146 </input>
<input>
<ID>IN_1</ID>147 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>166</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>61.5,-222.5</position>
<input>
<ID>IN_0</ID>162 </input>
<input>
<ID>IN_1</ID>163 </input>
<input>
<ID>IN_2</ID>164 </input>
<input>
<ID>IN_3</ID>165 </input>
<input>
<ID>IN_4</ID>166 </input>
<input>
<ID>IN_5</ID>167 </input>
<input>
<ID>IN_6</ID>168 </input>
<input>
<ID>IN_7</ID>169 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>165</ID>
<type>DD_KEYPAD_HEX</type>
<position>-63,-270.5</position>
<output>
<ID>OUT_0</ID>142 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>164</ID>
<type>AA_AND2</type>
<position>-31,-261.5</position>
<input>
<ID>IN_0</ID>138 </input>
<input>
<ID>IN_1</ID>139 </input>
<output>
<ID>OUT</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>162</ID>
<type>AI_XOR2</type>
<position>-17,-255.5</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>149 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>161</ID>
<type>AI_XOR2</type>
<position>19.5,-236.5</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>160 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>160</ID>
<type>AI_XOR2</type>
<position>-9.5,-261.5</position>
<input>
<ID>IN_0</ID>149 </input>
<input>
<ID>IN_1</ID>148 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_LABEL</type>
<position>-70.5,-270</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>AA_AND2</type>
<position>12,-225.5</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>157 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AI_XOR2</type>
<position>12,-230.5</position>
<input>
<ID>IN_0</ID>156 </input>
<input>
<ID>IN_1</ID>157 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>AA_AND2</type>
<position>-3,-236.5</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>152 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>155</ID>
<type>AA_AND2</type>
<position>4.5,-242.5</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>154 </input>
<output>
<ID>OUT</ID>153 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>154</ID>
<type>AE_OR2</type>
<position>10.5,-237.5</position>
<input>
<ID>IN_0</ID>152 </input>
<input>
<ID>IN_1</ID>153 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_AND2</type>
<position>-17,-250.5</position>
<input>
<ID>IN_0</ID>144 </input>
<input>
<ID>IN_1</ID>145 </input>
<output>
<ID>OUT</ID>146 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>152</ID>
<type>AE_OR2</type>
<position>25.5,-226.5</position>
<input>
<ID>IN_0</ID>158 </input>
<input>
<ID>IN_1</ID>159 </input>
<output>
<ID>OUT</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_AND2</type>
<position>19.5,-231.5</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>160 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>150</ID>
<type>AI_XOR2</type>
<position>4.5,-247.5</position>
<input>
<ID>IN_0</ID>155 </input>
<input>
<ID>IN_1</ID>154 </input>
<output>
<ID>OUT</ID>164 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>149</ID>
<type>AI_XOR2</type>
<position>-3,-241.5</position>
<input>
<ID>IN_0</ID>150 </input>
<input>
<ID>IN_1</ID>151 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>138</ID>
<type>AI_XOR2</type>
<position>-3,-189.5</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>119</ID>
<type>AI_XOR2</type>
<position>4.5,-195.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>168 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>AA_AND2</type>
<position>19.5,-179.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>136 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AE_OR2</type>
<position>25.5,-174.5</position>
<input>
<ID>IN_0</ID>134 </input>
<input>
<ID>IN_1</ID>135 </input>
<output>
<ID>OUT</ID>170 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_AND2</type>
<position>-17,-198.5</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>110</ID>
<type>AE_OR2</type>
<position>10.5,-185.5</position>
<input>
<ID>IN_0</ID>128 </input>
<input>
<ID>IN_1</ID>129 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>AA_AND2</type>
<position>4.5,-190.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>130 </input>
<output>
<ID>OUT</ID>129 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_AND2</type>
<position>-3,-184.5</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>127 </input>
<output>
<ID>OUT</ID>128 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>AI_XOR2</type>
<position>12,-178.5</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_AND2</type>
<position>12,-173.5</position>
<input>
<ID>IN_0</ID>132 </input>
<input>
<ID>IN_1</ID>133 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>105</ID>
<type>AI_XOR2</type>
<position>-9.5,-209.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>167 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AI_XOR2</type>
<position>19.5,-184.5</position>
<input>
<ID>IN_0</ID>137 </input>
<input>
<ID>IN_1</ID>136 </input>
<output>
<ID>OUT</ID>169 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>88</ID>
<type>AI_XOR2</type>
<position>-17,-203.5</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>-71,-190.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_AND2</type>
<position>-31,-209.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>66 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>-12.5,-168.5</position>
<gparam>LABEL_TEXT 8-Bits Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>DD_KEYPAD_HEX</type>
<position>-63,-190.5</position>
<output>
<ID>OUT_0</ID>32 </output>
<output>
<ID>OUT_1</ID>99 </output>
<output>
<ID>OUT_2</ID>126 </output>
<output>
<ID>OUT_3</ID>132 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>67</ID>
<type>AE_OR2</type>
<position>-3.5,-199.5</position>
<input>
<ID>IN_0</ID>113 </input>
<input>
<ID>IN_1</ID>114 </input>
<output>
<ID>OUT</ID>130 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>-71,-248</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_AND2</type>
<position>-23.5,-215.5</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>67 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>AI_XOR2</type>
<position>-31,-214.5</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>33 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>59</ID>
<type>AE_OR2</type>
<position>-17.5,-210.5</position>
<input>
<ID>IN_0</ID>66 </input>
<input>
<ID>IN_1</ID>67 </input>
<output>
<ID>OUT</ID>124 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AI_XOR2</type>
<position>-23.5,-220.5</position>
<input>
<ID>IN_0</ID>98 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>166 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_AND2</type>
<position>-9.5,-204.5</position>
<input>
<ID>IN_0</ID>125 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>114 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>DD_KEYPAD_HEX</type>
<position>-63,-235</position>
<output>
<ID>OUT_0</ID>33 </output>
<output>
<ID>OUT_1</ID>112 </output>
<output>
<ID>OUT_2</ID>127 </output>
<output>
<ID>OUT_3</ID>133 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>98</ID>
<type>DD_KEYPAD_HEX</type>
<position>69.5,5</position>
<output>
<ID>OUT_0</ID>25 </output>
<output>
<ID>OUT_1</ID>45 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 3</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>85,10.5</position>
<gparam>LABEL_TEXT 2-Bits Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>96</ID>
<type>DD_KEYPAD_HEX</type>
<position>69.5,-21</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>95</ID>
<type>AA_LABEL</type>
<position>62,-20.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_AND2</type>
<position>94,-8.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>93</ID>
<type>AI_XOR2</type>
<position>94,-13.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>92</ID>
<type>AE_OR2</type>
<position>100,-3.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>91</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>122,-12.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>51 </input>
<input>
<ID>IN_2</ID>52 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 5</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>90</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>45.5,-8</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 3</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>140</ID>
<type>AI_XOR2</type>
<position>-0.5,-63.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>DD_KEYPAD_HEX</type>
<position>69.5,-70</position>
<output>
<ID>OUT_0</ID>2 </output>
<output>
<ID>OUT_1</ID>10 </output>
<output>
<ID>OUT_2</ID>35 </output>
<output>
<ID>OUT_3</ID>41 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>81</ID>
<type>DD_KEYPAD_HEX</type>
<position>1,5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>139</ID>
<type>AI_XOR2</type>
<position>7,-69.5</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_AND2</type>
<position>108.5,-78</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>80</ID>
<type>DD_KEYPAD_HEX</type>
<position>1,-8</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_AND2</type>
<position>15.5,1</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>82</ID>
<type>AA_LABEL</type>
<position>16,11</position>
<gparam>LABEL_TEXT 1-Bit Full Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AA_AND2</type>
<position>22,-53.5</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AI_XOR2</type>
<position>94.5,-94</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>119 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>AE_OR2</type>
<position>28,-48.5</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>85 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AE_OR2</type>
<position>100.5,-84</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_AND2</type>
<position>-14.5,-72.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>65</ID>
<type>DD_KEYPAD_HEX</type>
<position>-46,5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>84</ID>
<type>DD_KEYPAD_HEX</type>
<position>1,-21</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>143</ID>
<type>AE_OR2</type>
<position>13,-59.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>AI_XOR2</type>
<position>87,-88</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>-6.5,-20.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND2</type>
<position>7,-64.5</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>17</ID>
<type>AA_AND2</type>
<position>94.5,-89</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>86</ID>
<type>AA_AND2</type>
<position>25.5,-7</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>145</ID>
<type>AA_AND2</type>
<position>-0.5,-58.5</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>62,-69.5</position>
<gparam>LABEL_TEXT B2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AI_XOR2</type>
<position>25.5,-14</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>21 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>146</ID>
<type>AI_XOR2</type>
<position>14.5,-52.5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>82 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>AE_OR2</type>
<position>114.5,-73</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>147</ID>
<type>AA_AND2</type>
<position>14.5,-47.5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>78 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>-31,11</position>
<gparam>LABEL_TEXT 1-Bit Half Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AI_XOR2</type>
<position>-7,-83.5</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>69 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>120</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>41,-73</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>69 </input>
<input>
<ID>IN_2</ID>83 </input>
<input>
<ID>IN_3</ID>84 </input>
<input>
<ID>IN_4</ID>85 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 15</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>121</ID>
<type>AE_OR2</type>
<position>-1,-73.5</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>63 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>-53.5,-70</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>AA_AND2</type>
<position>-21,-89.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>DD_KEYPAD_HEX</type>
<position>69.5,-57</position>
<output>
<ID>OUT_0</ID>1 </output>
<output>
<ID>OUT_1</ID>9 </output>
<output>
<ID>OUT_2</ID>34 </output>
<output>
<ID>OUT_3</ID>40 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>-6.5,5.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AI_XOR2</type>
<position>-28.5,-88.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>-37.5,17</position>
<gparam>LABEL_TEXT Logic Design HW2 412770116 </gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AE_OR2</type>
<position>114,7.5</position>
<input>
<ID>IN_0</ID>47 </input>
<input>
<ID>IN_1</ID>48 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>137</ID>
<type>AE_OR2</type>
<position>-15,-84.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>56 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>78</ID>
<type>AI_XOR2</type>
<position>15.5,-6</position>
<input>
<ID>IN_0</ID>13 </input>
<input>
<ID>IN_1</ID>14 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>AI_XOR2</type>
<position>-21,-94.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>68 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>105.5,-42</position>
<gparam>LABEL_TEXT 8-Bits Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>DD_KEYPAD_HEX</type>
<position>-46,-70.5</position>
<output>
<ID>OUT_0</ID>54 </output>
<output>
<ID>OUT_1</ID>61 </output>
<output>
<ID>OUT_2</ID>72 </output>
<output>
<ID>OUT_3</ID>78 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 7</lparam></gate>
<gate>
<ID>123</ID>
<type>AA_AND2</type>
<position>-7,-78.5</position>
<input>
<ID>IN_0</ID>65 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>134</ID>
<type>AA_LABEL</type>
<position>-53.5,-83</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_AND2</type>
<position>87,-83</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>-6.5,-7.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>133</ID>
<type>DD_KEYPAD_HEX</type>
<position>-46,-83.5</position>
<output>
<ID>OUT_0</ID>57 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>62,-56.5</position>
<gparam>LABEL_TEXT A2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>-53.5,-7.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>-10,-42.5</position>
<gparam>LABEL_TEXT 4-Bits Adder</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AI_XOR2</type>
<position>101,-77</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_LABEL</type>
<position>-53.5,5.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>72</ID>
<type>GE_LED_DISPLAY_4BIT</type>
<position>-20,-5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>11 </input>
<gparam>VALUE_BOX -1.9,-2.9,1.9,3.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 4</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>131</ID>
<type>DD_KEYPAD_HEX</type>
<position>-46,-57.5</position>
<output>
<ID>OUT_0</ID>53 </output>
<output>
<ID>OUT_1</ID>60 </output>
<output>
<ID>OUT_2</ID>71 </output>
<output>
<ID>OUT_3</ID>77 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 8</lparam></gate>
<gate>
<ID>4</ID>
<type>AI_XOR2</type>
<position>137.5,-58</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>122 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>AI_XOR2</type>
<position>-31.5,-6</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_AND2</type>
<position>-28.5,-83.5</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_AND2</type>
<position>-31.5,1</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>127</ID>
<type>AA_LABEL</type>
<position>-53.5,-57</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>AI_XOR2</type>
<position>-14.5,-77.5</position>
<input>
<ID>IN_0</ID>60 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>66</ID>
<type>DD_KEYPAD_HEX</type>
<position>-46,-8</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>89</ID>
<type>AE_OR2</type>
<position>35,0</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>AI_XOR2</type>
<position>22,-58.5</position>
<input>
<ID>IN_0</ID>82 </input>
<input>
<ID>IN_1</ID>81 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>21</ID>
<type>AI_XOR2</type>
<position>108.5,-83</position>
<input>
<ID>IN_0</ID>18 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>99</ID>
<type>DD_KEYPAD_HEX</type>
<position>69.5,-8</position>
<output>
<ID>OUT_0</ID>26 </output>
<output>
<ID>OUT_1</ID>46 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 2</lparam></gate>
<gate>
<ID>100</ID>
<type>AA_AND2</type>
<position>86.5,-2.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>101</ID>
<type>AI_XOR2</type>
<position>86.5,-7.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>102</ID>
<type>AA_LABEL</type>
<position>62,5.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>62,-7.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>AI_XOR2</type>
<position>100.5,3.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>AA_AND2</type>
<position>100.5,8.5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>46 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_AND2</type>
<position>108,2.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>117</ID>
<type>AI_XOR2</type>
<position>108,-2.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_AND2</type>
<position>130,-47</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>23</ID>
<type>AI_XOR2</type>
<position>130,-52</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_AND2</type>
<position>115,-58</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_AND2</type>
<position>122.5,-64</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>AE_OR2</type>
<position>128.5,-59</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>37 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>AA_AND2</type>
<position>101,-72</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AE_OR2</type>
<position>143.5,-48</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>123 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>AA_AND2</type>
<position>137.5,-53</position>
<input>
<ID>IN_0</ID>59 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AI_XOR2</type>
<position>122.5,-69</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>AI_XOR2</type>
<position>115,-63</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AI_XOR2</type>
<position>115,-115</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>33</ID>
<type>AI_XOR2</type>
<position>122.5,-121</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>117 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_AND2</type>
<position>137.5,-105</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>AE_OR2</type>
<position>143.5,-100</position>
<input>
<ID>IN_0</ID>108 </input>
<input>
<ID>IN_1</ID>109 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>AA_AND2</type>
<position>101,-124</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>AE_OR2</type>
<position>128.5,-111</position>
<input>
<ID>IN_0</ID>102 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_AND2</type>
<position>122.5,-116</position>
<input>
<ID>IN_0</ID>105 </input>
<input>
<ID>IN_1</ID>104 </input>
<output>
<ID>OUT</ID>103 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>AA_AND2</type>
<position>115,-110</position>
<input>
<ID>IN_0</ID>100 </input>
<input>
<ID>IN_1</ID>101 </input>
<output>
<ID>OUT</ID>102 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AI_XOR2</type>
<position>130,-104</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>41</ID>
<type>AA_AND2</type>
<position>130,-99</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>107 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>62,-134.5</position>
<gparam>LABEL_TEXT Carry</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AI_XOR2</type>
<position>108.5,-135</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>44</ID>
<type>AI_XOR2</type>
<position>137.5,-110</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>118 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>AI_XOR2</type>
<position>101,-129</position>
<input>
<ID>IN_0</ID>92 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>62,-108.5</position>
<gparam>LABEL_TEXT A1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_AND2</type>
<position>87,-135</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>48</ID>
<type>DD_KEYPAD_HEX</type>
<position>69.5,-135</position>
<output>
<ID>OUT_0</ID>90 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>50</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>179.5,-96</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>116 </input>
<input>
<ID>IN_2</ID>117 </input>
<input>
<ID>IN_3</ID>118 </input>
<input>
<ID>IN_4</ID>119 </input>
<input>
<ID>IN_5</ID>120 </input>
<input>
<ID>IN_6</ID>121 </input>
<input>
<ID>IN_7</ID>122 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 255</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>51</ID>
<type>AE_OR2</type>
<position>114.5,-125</position>
<input>
<ID>IN_0</ID>94 </input>
<input>
<ID>IN_1</ID>95 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>62,-121.5</position>
<gparam>LABEL_TEXT B1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_AND2</type>
<position>94.5,-141</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>AI_XOR2</type>
<position>87,-140</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>55</ID>
<type>AE_OR2</type>
<position>100.5,-136</position>
<input>
<ID>IN_0</ID>88 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>AI_XOR2</type>
<position>94.5,-146</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_AND2</type>
<position>108.5,-130</position>
<input>
<ID>IN_0</ID>97 </input>
<input>
<ID>IN_1</ID>96 </input>
<output>
<ID>OUT</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>DD_KEYPAD_HEX</type>
<position>69.5,-122</position>
<output>
<ID>OUT_0</ID>87 </output>
<output>
<ID>OUT_1</ID>93 </output>
<output>
<ID>OUT_2</ID>101 </output>
<output>
<ID>OUT_3</ID>107 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>49</ID>
<type>DD_KEYPAD_HEX</type>
<position>69.5,-109</position>
<output>
<ID>OUT_0</ID>86 </output>
<output>
<ID>OUT_1</ID>92 </output>
<output>
<ID>OUT_2</ID>100 </output>
<output>
<ID>OUT_3</ID>106 </output>
<gparam>KEYPAD_BOX_0 -3.65,3.05,-2.05,5.65</gparam>
<gparam>KEYPAD_BOX_1 -1.76,3.05,-0.16,5.65</gparam>
<gparam>KEYPAD_BOX_2 0.15,3.05,1.75,5.65</gparam>
<gparam>KEYPAD_BOX_3 2.05,3.05,3.65,5.65</gparam>
<gparam>KEYPAD_BOX_4 -3.65,0.15,-2.05,2.75</gparam>
<gparam>KEYPAD_BOX_5 -1.76,0.15,-0.16,2.75</gparam>
<gparam>KEYPAD_BOX_6 0.15,0.15,1.75,2.75</gparam>
<gparam>KEYPAD_BOX_7 2.05,0.15,3.65,2.75</gparam>
<gparam>KEYPAD_BOX_8 -3.65,-2.75,-2.05,-0.15</gparam>
<gparam>KEYPAD_BOX_9 -1.76,-2.75,-0.16,-0.15</gparam>
<gparam>KEYPAD_BOX_A 0.15,-2.75,1.75,-0.15</gparam>
<gparam>KEYPAD_BOX_B 2.05,-2.75,3.65,-0.15</gparam>
<gparam>KEYPAD_BOX_C -3.65,-5.65,-2.05,-3.05</gparam>
<gparam>KEYPAD_BOX_D -1.76,-5.65,-0.16,-3.05</gparam>
<gparam>KEYPAD_BOX_E 0.15,-5.65,1.75,-3.05</gparam>
<gparam>KEYPAD_BOX_F 2.05,-5.65,3.65,-3.05</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 4</lparam>
<lparam>OUTPUT_NUM 15</lparam></gate>
<gate>
<ID>60</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>179.5,-86.5</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<wire>
<ID>227 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320.5,-203.5,320.5,-162</points>
<intersection>-203.5 1</intersection>
<intersection>-162 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,-203.5,343,-203.5</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>320.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>315,-162,320.5,-162</points>
<connection>
<GID>210</GID>
<name>OUT</name></connection>
<intersection>320.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>226 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319.5,-206,319.5,-172</points>
<intersection>-206 1</intersection>
<intersection>-172 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319.5,-206,343,-206</points>
<connection>
<GID>190</GID>
<name>IN_7</name></connection>
<intersection>319.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309,-172,319.5,-172</points>
<connection>
<GID>218</GID>
<name>OUT</name></connection>
<intersection>319.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>225 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318.5,-207,318.5,-183</points>
<intersection>-207 1</intersection>
<intersection>-183 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318.5,-207,343,-207</points>
<connection>
<GID>190</GID>
<name>IN_6</name></connection>
<intersection>318.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>294,-183,318.5,-183</points>
<connection>
<GID>208</GID>
<name>OUT</name></connection>
<intersection>318.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>224 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317.5,-208,317.5,-197</points>
<intersection>-208 1</intersection>
<intersection>-197 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317.5,-208,343,-208</points>
<connection>
<GID>190</GID>
<name>IN_5</name></connection>
<intersection>317.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280,-197,317.5,-197</points>
<connection>
<GID>217</GID>
<name>OUT</name></connection>
<intersection>317.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>223 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>266,-209,343,-209</points>
<connection>
<GID>190</GID>
<name>IN_4</name></connection>
<intersection>266 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>266,-209,266,-208</points>
<connection>
<GID>229</GID>
<name>OUT</name></connection>
<intersection>-209 1</intersection></vsegment></shape></wire>
<wire>
<ID>222 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>317.5,-224,317.5,-210</points>
<intersection>-224 2</intersection>
<intersection>-210 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>317.5,-210,343,-210</points>
<connection>
<GID>190</GID>
<name>IN_3</name></connection>
<intersection>317.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>309,-224,317.5,-224</points>
<connection>
<GID>194</GID>
<name>OUT</name></connection>
<intersection>317.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>221 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>318.5,-235,318.5,-211</points>
<intersection>-235 2</intersection>
<intersection>-211 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>318.5,-211,343,-211</points>
<connection>
<GID>190</GID>
<name>IN_2</name></connection>
<intersection>318.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>294,-235,318.5,-235</points>
<connection>
<GID>205</GID>
<name>OUT</name></connection>
<intersection>318.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>220 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>319.5,-249,319.5,-212</points>
<intersection>-249 2</intersection>
<intersection>-212 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>319.5,-212,343,-212</points>
<connection>
<GID>190</GID>
<name>IN_1</name></connection>
<intersection>319.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>280,-249,319.5,-249</points>
<connection>
<GID>195</GID>
<name>OUT</name></connection>
<intersection>319.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>219 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>320.5,-260,320.5,-213</points>
<intersection>-260 2</intersection>
<intersection>-213 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>320.5,-213,343,-213</points>
<connection>
<GID>190</GID>
<name>IN_0</name></connection>
<intersection>320.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>266,-260,320.5,-260</points>
<connection>
<GID>185</GID>
<name>OUT</name></connection>
<intersection>320.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>218 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-223,301.5,-218</points>
<connection>
<GID>198</GID>
<name>OUT</name></connection>
<intersection>-223 23</intersection>
<intersection>-218 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-218,303,-218</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>301.5,-223,303,-223</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>217 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>300,-225,303,-225</points>
<connection>
<GID>201</GID>
<name>OUT</name></connection>
<connection>
<GID>194</GID>
<name>IN_1</name></connection>
<intersection>300 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>300,-225,300,-220</points>
<intersection>-225 1</intersection>
<intersection>-220 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>300,-220,303,-220</points>
<connection>
<GID>204</GID>
<name>IN_1</name></connection>
<intersection>300 3</intersection></hsegment></shape></wire>
<wire>
<ID>216 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-219,309,-215</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<connection>
<GID>204</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>215 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>301.5,-213,309,-213</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<connection>
<GID>197</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>214 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-219,294,-214</points>
<intersection>-219 2</intersection>
<intersection>-214 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>244.5,-219,295.5,-219</points>
<connection>
<GID>198</GID>
<name>IN_1</name></connection>
<intersection>244.5 8</intersection>
<intersection>294 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>244.5,-232.5,244.5,-219</points>
<intersection>-232.5 9</intersection>
<intersection>-219 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>228.5,-232.5,244.5,-232.5</points>
<connection>
<GID>183</GID>
<name>OUT_3</name></connection>
<intersection>244.5 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>294,-214,295.5,-214</points>
<connection>
<GID>197</GID>
<name>IN_1</name></connection>
<intersection>294 0</intersection></hsegment></shape></wire>
<wire>
<ID>213 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>292.5,-212,295.5,-212</points>
<connection>
<GID>197</GID>
<name>IN_0</name></connection>
<intersection>292.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>292.5,-217,292.5,-212</points>
<intersection>-217 4</intersection>
<intersection>-212 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>244,-217,295.5,-217</points>
<connection>
<GID>198</GID>
<name>IN_0</name></connection>
<intersection>244 9</intersection>
<intersection>292.5 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>244,-217,244,-188</points>
<intersection>-217 4</intersection>
<intersection>-188 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>228.5,-188,244,-188</points>
<connection>
<GID>182</GID>
<name>OUT_3</name></connection>
<intersection>244 9</intersection></hsegment></shape></wire>
<wire>
<ID>212 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>287,-234,287,-229</points>
<intersection>-234 23</intersection>
<intersection>-229 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>286.5,-229,288,-229</points>
<connection>
<GID>206</GID>
<name>OUT</name></connection>
<connection>
<GID>200</GID>
<name>IN_0</name></connection>
<intersection>287 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>287,-234,288,-234</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>287 0</intersection></hsegment></shape></wire>
<wire>
<ID>211 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>286,-236,288,-236</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>286 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>286,-239,286,-231</points>
<connection>
<GID>189</GID>
<name>OUT</name></connection>
<intersection>-236 1</intersection>
<intersection>-231 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>286,-231,288,-231</points>
<connection>
<GID>200</GID>
<name>IN_1</name></connection>
<intersection>286 12</intersection></hsegment></shape></wire>
<wire>
<ID>210 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-230,294,-226</points>
<connection>
<GID>200</GID>
<name>OUT</name></connection>
<connection>
<GID>201</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>209 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>286.5,-224,294,-224</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<connection>
<GID>199</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>208 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>278.5,-225,280.5,-225</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<intersection>278.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>278.5,-230,278.5,-225</points>
<intersection>-230 15</intersection>
<intersection>-225 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>245.5,-230,280.5,-230</points>
<connection>
<GID>206</GID>
<name>IN_1</name></connection>
<intersection>245.5 17</intersection>
<intersection>278.5 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>245.5,-234.5,245.5,-230</points>
<intersection>-234.5 18</intersection>
<intersection>-230 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>228.5,-234.5,245.5,-234.5</points>
<connection>
<GID>183</GID>
<name>OUT_2</name></connection>
<intersection>245.5 17</intersection></hsegment></shape></wire>
<wire>
<ID>207 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>245.5,-223,280.5,-223</points>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>245.5 20</intersection>
<intersection>276.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>276.5,-228,276.5,-223</points>
<intersection>-228 16</intersection>
<intersection>-223 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>276.5,-228,280.5,-228</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>276.5 12</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>245.5,-223,245.5,-190</points>
<intersection>-223 1</intersection>
<intersection>-190 27</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>228.5,-190,245.5,-190</points>
<connection>
<GID>182</GID>
<name>OUT_2</name></connection>
<intersection>245.5 20</intersection></hsegment></shape></wire>
<wire>
<ID>206 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>273,-248,273,-243</points>
<intersection>-248 23</intersection>
<intersection>-243 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>272.5,-243,274,-243</points>
<connection>
<GID>193</GID>
<name>OUT</name></connection>
<connection>
<GID>184</GID>
<name>IN_0</name></connection>
<intersection>273 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>273,-248,274,-248</points>
<connection>
<GID>195</GID>
<name>IN_0</name></connection>
<intersection>273 0</intersection></hsegment></shape></wire>
<wire>
<ID>205 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>272,-250,274,-250</points>
<connection>
<GID>195</GID>
<name>IN_1</name></connection>
<connection>
<GID>186</GID>
<name>OUT</name></connection>
<intersection>273.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>273.5,-250,273.5,-245</points>
<intersection>-250 1</intersection>
<intersection>-245 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>273.5,-245,274,-245</points>
<connection>
<GID>184</GID>
<name>IN_1</name></connection>
<intersection>273.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>204 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280,-244,280,-240</points>
<connection>
<GID>184</GID>
<name>OUT</name></connection>
<connection>
<GID>189</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>203 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>272.5,-238,280,-238</points>
<connection>
<GID>202</GID>
<name>OUT</name></connection>
<connection>
<GID>189</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>202 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,-244,264.5,-239</points>
<intersection>-244 2</intersection>
<intersection>-239 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>246,-244,266.5,-244</points>
<connection>
<GID>193</GID>
<name>IN_1</name></connection>
<intersection>246 8</intersection>
<intersection>264.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>264.5,-239,266.5,-239</points>
<connection>
<GID>202</GID>
<name>IN_1</name></connection>
<intersection>264.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>246,-244,246,-236.5</points>
<intersection>-244 2</intersection>
<intersection>-236.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>228.5,-236.5,246,-236.5</points>
<connection>
<GID>183</GID>
<name>OUT_1</name></connection>
<intersection>246 8</intersection></hsegment></shape></wire>
<wire>
<ID>201 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>246.5,-237,266.5,-237</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>246.5 6</intersection>
<intersection>263.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>263.5,-242,263.5,-237</points>
<intersection>-242 4</intersection>
<intersection>-237 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>263.5,-242,266.5,-242</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>263.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>246.5,-237,246.5,-192</points>
<intersection>-237 1</intersection>
<intersection>-192 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>228.5,-192,246.5,-192</points>
<connection>
<GID>182</GID>
<name>OUT_1</name></connection>
<intersection>246.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>200 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258.5,-259,258.5,-254</points>
<connection>
<GID>187</GID>
<name>OUT</name></connection>
<intersection>-259 23</intersection>
<intersection>-254 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>258.5,-254,260,-254</points>
<connection>
<GID>188</GID>
<name>IN_0</name></connection>
<intersection>258.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>258.5,-259,260,-259</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>258.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>199 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>228.5,-261,260,-261</points>
<connection>
<GID>191</GID>
<name>OUT_0</name></connection>
<connection>
<GID>185</GID>
<name>IN_1</name></connection>
<intersection>256.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>256.5,-261,256.5,-256</points>
<intersection>-261 1</intersection>
<intersection>-256 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>256.5,-256,260,-256</points>
<connection>
<GID>188</GID>
<name>IN_1</name></connection>
<intersection>256.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>198 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266,-255,266,-251</points>
<connection>
<GID>186</GID>
<name>IN_1</name></connection>
<connection>
<GID>188</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>197 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258.5,-249,266,-249</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>196 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>247,-250,252.5,-250</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<intersection>247 4</intersection>
<intersection>250 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>247,-250,247,-238.5</points>
<intersection>-250 2</intersection>
<intersection>-238.5 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>250,-255,250,-250</points>
<intersection>-255 15</intersection>
<intersection>-250 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>228.5,-238.5,247,-238.5</points>
<connection>
<GID>183</GID>
<name>OUT_0</name></connection>
<intersection>247 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>250,-255,252.5,-255</points>
<connection>
<GID>187</GID>
<name>IN_1</name></connection>
<intersection>250 11</intersection></hsegment></shape></wire>
<wire>
<ID>195 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>248,-248,252.5,-248</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>248 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>248,-253,248,-194</points>
<intersection>-253 16</intersection>
<intersection>-248 1</intersection>
<intersection>-194 24</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>248,-253,252.5,-253</points>
<connection>
<GID>187</GID>
<name>IN_0</name></connection>
<intersection>248 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>228.5,-194,248,-194</points>
<connection>
<GID>182</GID>
<name>OUT_0</name></connection>
<intersection>248 7</intersection></hsegment></shape></wire>
<wire>
<ID>194 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>301.5,-171,301.5,-166</points>
<connection>
<GID>215</GID>
<name>OUT</name></connection>
<intersection>-171 23</intersection>
<intersection>-166 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>301.5,-166,303,-166</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>301.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>301.5,-171,303,-171</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>301.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>193 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>300,-173,303,-173</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<connection>
<GID>212</GID>
<name>OUT</name></connection>
<intersection>301.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>301.5,-173,301.5,-168</points>
<intersection>-173 1</intersection>
<intersection>-168 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>301.5,-168,303,-168</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>301.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>192 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>309,-167,309,-163</points>
<connection>
<GID>209</GID>
<name>OUT</name></connection>
<connection>
<GID>210</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>191 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>301.5,-161,309,-161</points>
<connection>
<GID>216</GID>
<name>OUT</name></connection>
<connection>
<GID>210</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>190 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-167,294,-162</points>
<intersection>-167 2</intersection>
<intersection>-162 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>244.5,-167,295.5,-167</points>
<connection>
<GID>215</GID>
<name>IN_1</name></connection>
<intersection>244.5 8</intersection>
<intersection>294 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>244.5,-219.5,244.5,-167</points>
<intersection>-219.5 9</intersection>
<intersection>-167 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>228.5,-219.5,244.5,-219.5</points>
<connection>
<GID>231</GID>
<name>OUT_3</name></connection>
<intersection>244.5 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>294,-162,295.5,-162</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>294 0</intersection></hsegment></shape></wire>
<wire>
<ID>189 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>244,-160,295.5,-160</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>244 6</intersection>
<intersection>293 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>293,-165,293,-160</points>
<intersection>-165 4</intersection>
<intersection>-160 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>293,-165,295.5,-165</points>
<connection>
<GID>215</GID>
<name>IN_0</name></connection>
<intersection>293 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>244,-175,244,-160</points>
<intersection>-175 8</intersection>
<intersection>-160 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>228.5,-175,244,-175</points>
<connection>
<GID>223</GID>
<name>OUT_3</name></connection>
<intersection>244 6</intersection></hsegment></shape></wire>
<wire>
<ID>188 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>286.5,-182,286.5,-177</points>
<connection>
<GID>207</GID>
<name>OUT</name></connection>
<intersection>-182 23</intersection>
<intersection>-177 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>286.5,-177,288,-177</points>
<connection>
<GID>213</GID>
<name>IN_0</name></connection>
<intersection>286.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>286.5,-182,288,-182</points>
<connection>
<GID>208</GID>
<name>IN_0</name></connection>
<intersection>286.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>187 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>286,-184,288,-184</points>
<connection>
<GID>208</GID>
<name>IN_1</name></connection>
<intersection>286 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>286,-187,286,-179</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<intersection>-184 1</intersection>
<intersection>-179 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>286,-179,288,-179</points>
<connection>
<GID>213</GID>
<name>IN_1</name></connection>
<intersection>286 12</intersection></hsegment></shape></wire>
<wire>
<ID>186 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>294,-178,294,-174</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<connection>
<GID>213</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>185 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>286.5,-172,294,-172</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<connection>
<GID>212</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>184 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>278.5,-173,280.5,-173</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>278.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>278.5,-178,278.5,-173</points>
<intersection>-178 15</intersection>
<intersection>-173 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>245,-178,280.5,-178</points>
<connection>
<GID>207</GID>
<name>IN_1</name></connection>
<intersection>245 17</intersection>
<intersection>278.5 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>245,-221.5,245,-178</points>
<intersection>-221.5 18</intersection>
<intersection>-178 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>228.5,-221.5,245,-221.5</points>
<connection>
<GID>231</GID>
<name>OUT_2</name></connection>
<intersection>245 17</intersection></hsegment></shape></wire>
<wire>
<ID>183 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>228.5,-177,280.5,-177</points>
<connection>
<GID>223</GID>
<name>OUT_2</name></connection>
<intersection>275.5 20</intersection>
<intersection>280.5 23</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>275.5,-177,275.5,-171</points>
<intersection>-177 1</intersection>
<intersection>-171 22</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>275.5,-171,280.5,-171</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>275.5 20</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>280.5,-177,280.5,-176</points>
<connection>
<GID>207</GID>
<name>IN_0</name></connection>
<intersection>-177 1</intersection></vsegment></shape></wire>
<wire>
<ID>182 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>272.5,-196,272.5,-191</points>
<connection>
<GID>219</GID>
<name>OUT</name></connection>
<intersection>-196 23</intersection>
<intersection>-191 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>272.5,-191,274,-191</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>272.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>272.5,-196,274,-196</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<intersection>272.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>181 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>272,-198,274,-198</points>
<connection>
<GID>217</GID>
<name>IN_1</name></connection>
<intersection>272 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>272,-198,272,-193</points>
<connection>
<GID>228</GID>
<name>OUT</name></connection>
<intersection>-198 1</intersection>
<intersection>-193 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>272,-193,274,-193</points>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<intersection>272 3</intersection></hsegment></shape></wire>
<wire>
<ID>180 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>280,-192,280,-188</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<connection>
<GID>230</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>179 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>272.5,-186,280,-186</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<connection>
<GID>211</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>178 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>264.5,-192,264.5,-187</points>
<intersection>-192 2</intersection>
<intersection>-187 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>246,-192,266.5,-192</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>246 8</intersection>
<intersection>264.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>264.5,-187,266.5,-187</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<intersection>264.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>246,-223.5,246,-192</points>
<intersection>-223.5 9</intersection>
<intersection>-192 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>228.5,-223.5,246,-223.5</points>
<connection>
<GID>231</GID>
<name>OUT_1</name></connection>
<intersection>246 8</intersection></hsegment></shape></wire>
<wire>
<ID>177 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>228.5,-179,266.5,-179</points>
<connection>
<GID>223</GID>
<name>OUT_1</name></connection>
<intersection>266.5 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>266.5,-190,266.5,-179</points>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>-179 1</intersection></vsegment></shape></wire>
<wire>
<ID>176 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>258.5,-207,258.5,-202</points>
<connection>
<GID>227</GID>
<name>OUT</name></connection>
<intersection>-207 23</intersection>
<intersection>-202 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>258.5,-202,260,-202</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>258.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>258.5,-207,260,-207</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>258.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>175 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>256.5,-210.5,316.5,-210.5</points>
<intersection>256.5 12</intersection>
<intersection>260 19</intersection>
<intersection>316.5 15</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>256.5,-210.5,256.5,-204</points>
<intersection>-210.5 1</intersection>
<intersection>-204 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>256.5,-204,260,-204</points>
<connection>
<GID>226</GID>
<name>IN_1</name></connection>
<intersection>256.5 12</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>316.5,-214,316.5,-210.5</points>
<intersection>-214 32</intersection>
<intersection>-210.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>260,-210.5,260,-209</points>
<connection>
<GID>229</GID>
<name>IN_1</name></connection>
<intersection>-210.5 1</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>315,-214,316.5,-214</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>316.5 15</intersection></hsegment></shape></wire>
<wire>
<ID>174 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>266,-203,266,-199</points>
<connection>
<GID>226</GID>
<name>OUT</name></connection>
<connection>
<GID>228</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>173 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>258.5,-197,266,-197</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<connection>
<GID>221</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>172 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>247,-198,252.5,-198</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>247 4</intersection>
<intersection>250 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>247,-225.5,247,-198</points>
<intersection>-225.5 14</intersection>
<intersection>-198 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>250,-203,250,-198</points>
<intersection>-203 15</intersection>
<intersection>-198 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>228.5,-225.5,247,-225.5</points>
<connection>
<GID>231</GID>
<name>OUT_0</name></connection>
<intersection>247 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>250,-203,252.5,-203</points>
<connection>
<GID>227</GID>
<name>IN_1</name></connection>
<intersection>250 11</intersection></hsegment></shape></wire>
<wire>
<ID>171 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>248,-196,252.5,-196</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>248 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>248,-201,248,-181</points>
<intersection>-201 16</intersection>
<intersection>-196 1</intersection>
<intersection>-181 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>228.5,-181,248,-181</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>248 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>248,-201,252.5,-201</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>248 7</intersection></hsegment></shape></wire>
<wire>
<ID>170 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-216,34,-174.5</points>
<intersection>-216 1</intersection>
<intersection>-174.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-216,56.5,-216</points>
<connection>
<GID>176</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-174.5,34,-174.5</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>169 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-218.5,33,-184.5</points>
<intersection>-218.5 1</intersection>
<intersection>-184.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-218.5,56.5,-218.5</points>
<connection>
<GID>166</GID>
<name>IN_7</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-184.5,33,-184.5</points>
<connection>
<GID>104</GID>
<name>OUT</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>168 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-219.5,32,-195.5</points>
<intersection>-219.5 1</intersection>
<intersection>-195.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-219.5,56.5,-219.5</points>
<connection>
<GID>166</GID>
<name>IN_6</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-195.5,32,-195.5</points>
<connection>
<GID>119</GID>
<name>OUT</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>167 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-220.5,31,-209.5</points>
<intersection>-220.5 1</intersection>
<intersection>-209.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-220.5,56.5,-220.5</points>
<connection>
<GID>166</GID>
<name>IN_5</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6.5,-209.5,31,-209.5</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>166 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20.5,-221.5,56.5,-221.5</points>
<connection>
<GID>166</GID>
<name>IN_4</name></connection>
<intersection>-20.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-20.5,-221.5,-20.5,-220.5</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<intersection>-221.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>165 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-236.5,31,-222.5</points>
<intersection>-236.5 2</intersection>
<intersection>-222.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-222.5,56.5,-222.5</points>
<connection>
<GID>166</GID>
<name>IN_3</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>22.5,-236.5,31,-236.5</points>
<connection>
<GID>161</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>164 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>32,-247.5,32,-223.5</points>
<intersection>-247.5 2</intersection>
<intersection>-223.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-223.5,56.5,-223.5</points>
<connection>
<GID>166</GID>
<name>IN_2</name></connection>
<intersection>32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>7.5,-247.5,32,-247.5</points>
<connection>
<GID>150</GID>
<name>OUT</name></connection>
<intersection>32 0</intersection></hsegment></shape></wire>
<wire>
<ID>163 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-261.5,33,-224.5</points>
<intersection>-261.5 2</intersection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-224.5,56.5,-224.5</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6.5,-261.5,33,-261.5</points>
<connection>
<GID>160</GID>
<name>OUT</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>162 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-272.5,34,-225.5</points>
<intersection>-272.5 2</intersection>
<intersection>-225.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>34,-225.5,56.5,-225.5</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-20.5,-272.5,34,-272.5</points>
<connection>
<GID>172</GID>
<name>OUT</name></connection>
<intersection>34 0</intersection></hsegment></shape></wire>
<wire>
<ID>161 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-235.5,15,-230.5</points>
<connection>
<GID>157</GID>
<name>OUT</name></connection>
<intersection>-235.5 23</intersection>
<intersection>-230.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>15,-230.5,16.5,-230.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>15,-235.5,16.5,-235.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>160 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-237.5,16.5,-237.5</points>
<connection>
<GID>161</GID>
<name>IN_1</name></connection>
<connection>
<GID>154</GID>
<name>OUT</name></connection>
<intersection>13.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13.5,-237.5,13.5,-232.5</points>
<intersection>-237.5 1</intersection>
<intersection>-232.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>13.5,-232.5,16.5,-232.5</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<intersection>13.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>159 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-231.5,22.5,-227.5</points>
<connection>
<GID>151</GID>
<name>OUT</name></connection>
<connection>
<GID>152</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>158 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-225.5,22.5,-225.5</points>
<connection>
<GID>158</GID>
<name>OUT</name></connection>
<connection>
<GID>152</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>157 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-231.5,7.5,-226.5</points>
<intersection>-231.5 2</intersection>
<intersection>-226.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-42,-231.5,9,-231.5</points>
<connection>
<GID>157</GID>
<name>IN_1</name></connection>
<intersection>-42 8</intersection>
<intersection>7.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-42,-245,-42,-231.5</points>
<intersection>-245 9</intersection>
<intersection>-231.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-58,-245,-42,-245</points>
<connection>
<GID>174</GID>
<name>OUT_3</name></connection>
<intersection>-42 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>7.5,-226.5,9,-226.5</points>
<connection>
<GID>158</GID>
<name>IN_1</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>156 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,-224.5,9,-224.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>6 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>6,-229.5,6,-224.5</points>
<intersection>-229.5 4</intersection>
<intersection>-224.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-42.5,-229.5,9,-229.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>-42.5 9</intersection>
<intersection>6 3</intersection></hsegment>
<vsegment>
<ID>9</ID>
<points>-42.5,-229.5,-42.5,-200.5</points>
<intersection>-229.5 4</intersection>
<intersection>-200.5 10</intersection></vsegment>
<hsegment>
<ID>10</ID>
<points>-58,-200.5,-42.5,-200.5</points>
<connection>
<GID>175</GID>
<name>OUT_3</name></connection>
<intersection>-42.5 9</intersection></hsegment></shape></wire>
<wire>
<ID>155 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0.5,-246.5,0.5,-241.5</points>
<intersection>-246.5 23</intersection>
<intersection>-241.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>0,-241.5,1.5,-241.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>0.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>0.5,-246.5,1.5,-246.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>0.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>154 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-248.5,1.5,-248.5</points>
<connection>
<GID>150</GID>
<name>IN_1</name></connection>
<intersection>-0.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-0.5,-251.5,-0.5,-243.5</points>
<connection>
<GID>167</GID>
<name>OUT</name></connection>
<intersection>-248.5 1</intersection>
<intersection>-243.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-0.5,-243.5,1.5,-243.5</points>
<connection>
<GID>155</GID>
<name>IN_1</name></connection>
<intersection>-0.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>153 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-242.5,7.5,-238.5</points>
<connection>
<GID>154</GID>
<name>IN_1</name></connection>
<connection>
<GID>155</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>152 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-236.5,7.5,-236.5</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<connection>
<GID>154</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>151 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-8,-237.5,-6,-237.5</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>-8 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-8,-242.5,-8,-237.5</points>
<intersection>-242.5 15</intersection>
<intersection>-237.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-41,-242.5,-6,-242.5</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>-41 17</intersection>
<intersection>-8 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>-41,-247,-41,-242.5</points>
<intersection>-247 18</intersection>
<intersection>-242.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-58,-247,-41,-247</points>
<connection>
<GID>174</GID>
<name>OUT_2</name></connection>
<intersection>-41 17</intersection></hsegment></shape></wire>
<wire>
<ID>150 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-235.5,-6,-235.5</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>-41 20</intersection>
<intersection>-10 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-10,-240.5,-10,-235.5</points>
<intersection>-240.5 16</intersection>
<intersection>-235.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-10,-240.5,-6,-240.5</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>-10 12</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>-41,-235.5,-41,-202.5</points>
<intersection>-235.5 1</intersection>
<intersection>-202.5 27</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>-58,-202.5,-41,-202.5</points>
<connection>
<GID>175</GID>
<name>OUT_2</name></connection>
<intersection>-41 20</intersection></hsegment></shape></wire>
<wire>
<ID>149 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-13.5,-260.5,-13.5,-255.5</points>
<intersection>-260.5 23</intersection>
<intersection>-255.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14,-255.5,-12.5,-255.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<connection>
<GID>162</GID>
<name>OUT</name></connection>
<intersection>-13.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-13.5,-260.5,-12.5,-260.5</points>
<connection>
<GID>160</GID>
<name>IN_0</name></connection>
<intersection>-13.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>148 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14.5,-262.5,-12.5,-262.5</points>
<connection>
<GID>171</GID>
<name>OUT</name></connection>
<connection>
<GID>160</GID>
<name>IN_1</name></connection>
<intersection>-14.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-14.5,-262.5,-14.5,-257.5</points>
<intersection>-262.5 1</intersection>
<intersection>-257.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-14.5,-257.5,-12.5,-257.5</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>-14.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>147 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,-256.5,-6.5,-252.5</points>
<connection>
<GID>167</GID>
<name>IN_1</name></connection>
<connection>
<GID>173</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>146 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14,-250.5,-6.5,-250.5</points>
<connection>
<GID>153</GID>
<name>OUT</name></connection>
<connection>
<GID>167</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>145 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-256.5,-22,-251.5</points>
<intersection>-256.5 2</intersection>
<intersection>-251.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-40.5,-256.5,-20,-256.5</points>
<connection>
<GID>162</GID>
<name>IN_1</name></connection>
<intersection>-40.5 8</intersection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-22,-251.5,-20,-251.5</points>
<connection>
<GID>153</GID>
<name>IN_1</name></connection>
<intersection>-22 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-40.5,-256.5,-40.5,-249</points>
<intersection>-256.5 2</intersection>
<intersection>-249 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-58,-249,-40.5,-249</points>
<connection>
<GID>174</GID>
<name>OUT_1</name></connection>
<intersection>-40.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>144 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-249.5,-20,-249.5</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>-40 6</intersection>
<intersection>-23 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-23,-254.5,-23,-249.5</points>
<intersection>-254.5 4</intersection>
<intersection>-249.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-23,-254.5,-20,-254.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>-23 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-40,-249.5,-40,-204.5</points>
<intersection>-249.5 1</intersection>
<intersection>-204.5 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>-58,-204.5,-40,-204.5</points>
<connection>
<GID>175</GID>
<name>OUT_1</name></connection>
<intersection>-40 6</intersection></hsegment></shape></wire>
<wire>
<ID>143 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-271.5,-28,-266.5</points>
<connection>
<GID>170</GID>
<name>OUT</name></connection>
<intersection>-271.5 23</intersection>
<intersection>-266.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-28,-266.5,-26.5,-266.5</points>
<connection>
<GID>169</GID>
<name>IN_0</name></connection>
<intersection>-28 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-28,-271.5,-26.5,-271.5</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>-28 0</intersection></hsegment></shape></wire>
<wire>
<ID>142 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-58,-273.5,-26.5,-273.5</points>
<connection>
<GID>172</GID>
<name>IN_1</name></connection>
<connection>
<GID>165</GID>
<name>OUT_0</name></connection>
<intersection>-30 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-30,-273.5,-30,-268.5</points>
<intersection>-273.5 1</intersection>
<intersection>-268.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-30,-268.5,-26.5,-268.5</points>
<connection>
<GID>169</GID>
<name>IN_1</name></connection>
<intersection>-30 12</intersection></hsegment></shape></wire>
<wire>
<ID>141 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,-267.5,-20.5,-263.5</points>
<connection>
<GID>169</GID>
<name>OUT</name></connection>
<connection>
<GID>171</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>140 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28,-261.5,-20.5,-261.5</points>
<connection>
<GID>164</GID>
<name>OUT</name></connection>
<connection>
<GID>171</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>139 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-39.5,-262.5,-34,-262.5</points>
<connection>
<GID>164</GID>
<name>IN_1</name></connection>
<intersection>-39.5 4</intersection>
<intersection>-36.5 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-39.5,-262.5,-39.5,-251</points>
<intersection>-262.5 2</intersection>
<intersection>-251 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-36.5,-267.5,-36.5,-262.5</points>
<intersection>-267.5 15</intersection>
<intersection>-262.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-58,-251,-39.5,-251</points>
<connection>
<GID>174</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-36.5,-267.5,-34,-267.5</points>
<connection>
<GID>170</GID>
<name>IN_1</name></connection>
<intersection>-36.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>138 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-38.5,-260.5,-34,-260.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>-38.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-38.5,-265.5,-38.5,-206.5</points>
<intersection>-265.5 16</intersection>
<intersection>-260.5 1</intersection>
<intersection>-206.5 24</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-38.5,-265.5,-34,-265.5</points>
<connection>
<GID>170</GID>
<name>IN_0</name></connection>
<intersection>-38.5 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>-58,-206.5,-38.5,-206.5</points>
<connection>
<GID>175</GID>
<name>OUT_0</name></connection>
<intersection>-38.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>137 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15,-183.5,15,-178.5</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<intersection>-183.5 23</intersection>
<intersection>-178.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>15,-178.5,16.5,-178.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>15,-183.5,16.5,-183.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>15 0</intersection></hsegment></shape></wire>
<wire>
<ID>136 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-185.5,16.5,-185.5</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<intersection>13.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>13.5,-185.5,13.5,-180.5</points>
<intersection>-185.5 1</intersection>
<intersection>-180.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>13.5,-180.5,16.5,-180.5</points>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>13.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>135 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>22.5,-179.5,22.5,-175.5</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<connection>
<GID>113</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>134 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>15,-173.5,22.5,-173.5</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<connection>
<GID>112</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>133 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-179.5,7.5,-174.5</points>
<intersection>-179.5 2</intersection>
<intersection>-174.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-42,-179.5,9,-179.5</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>-42 8</intersection>
<intersection>7.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-42,-232,-42,-179.5</points>
<intersection>-232 9</intersection>
<intersection>-179.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-58,-232,-42,-232</points>
<connection>
<GID>10</GID>
<name>OUT_3</name></connection>
<intersection>-42 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>7.5,-174.5,9,-174.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>7.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-42.5,-172.5,9,-172.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>-42.5 6</intersection>
<intersection>6.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>6.5,-177.5,6.5,-172.5</points>
<intersection>-177.5 4</intersection>
<intersection>-172.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>6.5,-177.5,9,-177.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>6.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-42.5,-187.5,-42.5,-172.5</points>
<intersection>-187.5 8</intersection>
<intersection>-172.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-58,-187.5,-42.5,-187.5</points>
<connection>
<GID>69</GID>
<name>OUT_3</name></connection>
<intersection>-42.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>131 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>0,-194.5,0,-189.5</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>-194.5 23</intersection>
<intersection>-189.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>0,-189.5,1.5,-189.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>0 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>0,-194.5,1.5,-194.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>0 0</intersection></hsegment></shape></wire>
<wire>
<ID>130 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-0.5,-196.5,1.5,-196.5</points>
<connection>
<GID>119</GID>
<name>IN_1</name></connection>
<intersection>-0.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-0.5,-199.5,-0.5,-191.5</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>-196.5 1</intersection>
<intersection>-191.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-0.5,-191.5,1.5,-191.5</points>
<connection>
<GID>109</GID>
<name>IN_1</name></connection>
<intersection>-0.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>129 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>7.5,-190.5,7.5,-186.5</points>
<connection>
<GID>109</GID>
<name>OUT</name></connection>
<connection>
<GID>110</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>128 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>0,-184.5,7.5,-184.5</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<connection>
<GID>110</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>127 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-8,-185.5,-6,-185.5</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>-8 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-8,-190.5,-8,-185.5</points>
<intersection>-190.5 15</intersection>
<intersection>-185.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-41.5,-190.5,-6,-190.5</points>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>-41.5 17</intersection>
<intersection>-8 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>-41.5,-234,-41.5,-190.5</points>
<intersection>-234 18</intersection>
<intersection>-190.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-58,-234,-41.5,-234</points>
<connection>
<GID>10</GID>
<name>OUT_2</name></connection>
<intersection>-41.5 17</intersection></hsegment></shape></wire>
<wire>
<ID>126 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-58,-189.5,-6,-189.5</points>
<connection>
<GID>69</GID>
<name>OUT_2</name></connection>
<intersection>-11 20</intersection>
<intersection>-6 23</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>-11,-189.5,-11,-183.5</points>
<intersection>-189.5 1</intersection>
<intersection>-183.5 22</intersection></vsegment>
<hsegment>
<ID>22</ID>
<points>-11,-183.5,-6,-183.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>-11 20</intersection></hsegment>
<vsegment>
<ID>23</ID>
<points>-6,-189.5,-6,-188.5</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>-189.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>125 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-14,-208.5,-14,-203.5</points>
<connection>
<GID>88</GID>
<name>OUT</name></connection>
<intersection>-208.5 23</intersection>
<intersection>-203.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-14,-203.5,-12.5,-203.5</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-14,-208.5,-12.5,-208.5</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>-14 0</intersection></hsegment></shape></wire>
<wire>
<ID>124 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14.5,-210.5,-12.5,-210.5</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<intersection>-14.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-14.5,-210.5,-14.5,-205.5</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<intersection>-210.5 1</intersection>
<intersection>-205.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-14.5,-205.5,-12.5,-205.5</points>
<connection>
<GID>11</GID>
<name>IN_1</name></connection>
<intersection>-14.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>114 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-6.5,-204.5,-6.5,-200.5</points>
<connection>
<GID>11</GID>
<name>OUT</name></connection>
<connection>
<GID>67</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>113 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14,-198.5,-6.5,-198.5</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<connection>
<GID>67</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>112 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-22,-204.5,-22,-199.5</points>
<intersection>-204.5 2</intersection>
<intersection>-199.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-40.5,-204.5,-20,-204.5</points>
<connection>
<GID>88</GID>
<name>IN_1</name></connection>
<intersection>-40.5 8</intersection>
<intersection>-22 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-22,-199.5,-20,-199.5</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>-22 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-40.5,-236,-40.5,-204.5</points>
<intersection>-236 9</intersection>
<intersection>-204.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-58,-236,-40.5,-236</points>
<connection>
<GID>10</GID>
<name>OUT_1</name></connection>
<intersection>-40.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>99 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-58,-191.5,-20,-191.5</points>
<connection>
<GID>69</GID>
<name>OUT_1</name></connection>
<intersection>-20 6</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-20,-202.5,-20,-191.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<connection>
<GID>88</GID>
<name>IN_0</name></connection>
<intersection>-191.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>98 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-28,-219.5,-28,-214.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>-219.5 23</intersection>
<intersection>-214.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-28,-214.5,-26.5,-214.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-28 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-28,-219.5,-26.5,-219.5</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>-28 0</intersection></hsegment></shape></wire>
<wire>
<ID>70 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-30,-223,30,-223</points>
<intersection>-30 12</intersection>
<intersection>-26.5 19</intersection>
<intersection>30 15</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-30,-223,-30,-216.5</points>
<intersection>-223 1</intersection>
<intersection>-216.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-30,-216.5,-26.5,-216.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>-30 12</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>30,-226.5,30,-223</points>
<intersection>-226.5 32</intersection>
<intersection>-223 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>-26.5,-223,-26.5,-221.5</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<intersection>-223 1</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>28.5,-226.5,30,-226.5</points>
<connection>
<GID>152</GID>
<name>OUT</name></connection>
<intersection>30 15</intersection></hsegment></shape></wire>
<wire>
<ID>67 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,-215.5,-20.5,-211.5</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<connection>
<GID>62</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>66 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28,-209.5,-20.5,-209.5</points>
<connection>
<GID>77</GID>
<name>OUT</name></connection>
<connection>
<GID>59</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-39.5,-210.5,-34,-210.5</points>
<connection>
<GID>77</GID>
<name>IN_1</name></connection>
<intersection>-39.5 4</intersection>
<intersection>-36.5 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-39.5,-238,-39.5,-210.5</points>
<intersection>-238 14</intersection>
<intersection>-210.5 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-36.5,-215.5,-36.5,-210.5</points>
<intersection>-215.5 15</intersection>
<intersection>-210.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-58,-238,-39.5,-238</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-39.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-36.5,-215.5,-34,-215.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>-36.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>32 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-38.5,-208.5,-34,-208.5</points>
<connection>
<GID>77</GID>
<name>IN_0</name></connection>
<intersection>-38.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-38.5,-213.5,-38.5,-193.5</points>
<intersection>-213.5 16</intersection>
<intersection>-208.5 1</intersection>
<intersection>-193.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-58,-193.5,-38.5,-193.5</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>-38.5 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-38.5,-213.5,-34,-213.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>-38.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>29 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>82,-24,82,-14.5</points>
<intersection>-24 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82,-14.5,91,-14.5</points>
<connection>
<GID>93</GID>
<name>IN_1</name></connection>
<intersection>82 0</intersection>
<intersection>85.5 12</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74.5,-24,82,-24</points>
<connection>
<GID>96</GID>
<name>OUT_0</name></connection>
<intersection>82 0</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>85.5,-14.5,85.5,-9.5</points>
<intersection>-14.5 1</intersection>
<intersection>-9.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>85.5,-9.5,91,-9.5</points>
<connection>
<GID>94</GID>
<name>IN_1</name></connection>
<intersection>85.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>28 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97,-8.5,97,-4.5</points>
<connection>
<GID>92</GID>
<name>IN_1</name></connection>
<connection>
<GID>94</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>31 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,-13.5,119,-13.5</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<connection>
<GID>93</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>80 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>25,-53.5,25,-49.5</points>
<connection>
<GID>141</GID>
<name>OUT</name></connection>
<connection>
<GID>142</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>74 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-64.5,10,-60.5</points>
<connection>
<GID>143</GID>
<name>IN_1</name></connection>
<connection>
<GID>144</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>76 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2.5,-68.5,2.5,-63.5</points>
<connection>
<GID>140</GID>
<name>OUT</name></connection>
<intersection>-68.5 23</intersection>
<intersection>-63.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>2.5,-63.5,4,-63.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>2.5,-68.5,4,-68.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-89,97.5,-85</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<connection>
<GID>17</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>8 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-93,90,-88</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>-93 23</intersection>
<intersection>-88 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>90,-88,91.5,-88</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>90,-93,91.5,-93</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>73 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2.5,-58.5,10,-58.5</points>
<connection>
<GID>143</GID>
<name>IN_0</name></connection>
<connection>
<GID>145</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>23 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-14,39.5,-9</points>
<intersection>-14 2</intersection>
<intersection>-9 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-9,42.5,-9</points>
<connection>
<GID>90</GID>
<name>IN_0</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-14,39.5,-14</points>
<connection>
<GID>87</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13.5,-24,13.5,-15</points>
<intersection>-24 2</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>13.5,-15,22.5,-15</points>
<connection>
<GID>87</GID>
<name>IN_1</name></connection>
<intersection>13.5 0</intersection>
<intersection>19 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-24,13.5,-24</points>
<connection>
<GID>84</GID>
<name>OUT_0</name></connection>
<intersection>13.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>19,-15,19,-8</points>
<intersection>-15 1</intersection>
<intersection>-8 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>19,-8,22.5,-8</points>
<connection>
<GID>86</GID>
<name>IN_1</name></connection>
<intersection>19 3</intersection></hsegment></shape></wire>
<wire>
<ID>16 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-78,111.5,-74</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>19</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>79 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>17.5,-47.5,25,-47.5</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<connection>
<GID>147</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>85 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-72,35,-48.5</points>
<intersection>-72 1</intersection>
<intersection>-48.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>35,-72,36,-72</points>
<connection>
<GID>120</GID>
<name>IN_4</name></connection>
<intersection>35 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-48.5,35,-48.5</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>83 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>15.5,-74,15.5,-69.5</points>
<intersection>-74 1</intersection>
<intersection>-69.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>15.5,-74,36,-74</points>
<connection>
<GID>120</GID>
<name>IN_2</name></connection>
<intersection>15.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>10,-69.5,15.5,-69.5</points>
<connection>
<GID>139</GID>
<name>OUT</name></connection>
<intersection>15.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>8.5,-83.5,8.5,-75</points>
<intersection>-83.5 2</intersection>
<intersection>-75 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>8.5,-75,36,-75</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>8.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-4,-83.5,8.5,-83.5</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>8.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>2,-70.5,4,-70.5</points>
<connection>
<GID>139</GID>
<name>IN_1</name></connection>
<intersection>2 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>2,-73.5,2,-65.5</points>
<connection>
<GID>121</GID>
<name>OUT</name></connection>
<intersection>-70.5 1</intersection>
<intersection>-65.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>2,-65.5,4,-65.5</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>2 12</intersection></hsegment></shape></wire>
<wire>
<ID>62 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-11.5,-72.5,-4,-72.5</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<connection>
<GID>124</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>52 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-11.5,118,7.5</points>
<intersection>-11.5 1</intersection>
<intersection>7.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>118,-11.5,119,-11.5</points>
<connection>
<GID>91</GID>
<name>IN_2</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>117,7.5,118,7.5</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>56 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-18,-89.5,-18,-85.5</points>
<connection>
<GID>137</GID>
<name>IN_1</name></connection>
<connection>
<GID>135</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>22 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-13,20.5,-6</points>
<intersection>-13 1</intersection>
<intersection>-6 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-13,22.5,-13</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>18.5,-6,22.5,-6</points>
<connection>
<GID>78</GID>
<name>OUT</name></connection>
<connection>
<GID>86</GID>
<name>IN_0</name></connection>
<intersection>20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-11,10,0</points>
<intersection>-11 2</intersection>
<intersection>-7 3</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,0,12.5,0</points>
<connection>
<GID>79</GID>
<name>IN_1</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>6,-11,10,-11</points>
<connection>
<GID>80</GID>
<name>OUT_0</name></connection>
<intersection>10 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>10,-7,12.5,-7</points>
<connection>
<GID>78</GID>
<name>IN_1</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>13 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>6,2,12.5,2</points>
<connection>
<GID>81</GID>
<name>OUT_0</name></connection>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>8 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>8,-5,8,2</points>
<intersection>-5 4</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>8,-5,12.5,-5</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>8 3</intersection></hsegment></shape></wire>
<wire>
<ID>68 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18,-94.5,35,-94.5</points>
<connection>
<GID>136</GID>
<name>OUT</name></connection>
<intersection>35 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>35,-94.5,35,-76</points>
<intersection>-94.5 1</intersection>
<intersection>-76 12</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>35,-76,36,-76</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>35 11</intersection></hsegment></shape></wire>
<wire>
<ID>58 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,-93.5,-25.5,-88.5</points>
<connection>
<GID>128</GID>
<name>OUT</name></connection>
<intersection>-93.5 23</intersection>
<intersection>-88.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-25.5,-88.5,-24,-88.5</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-25.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-25.5,-93.5,-24,-93.5</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>-25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>78 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>10,-53.5,10,-48.5</points>
<intersection>-53.5 2</intersection>
<intersection>-48.5 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-39.5,-53.5,11.5,-53.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>-39.5 8</intersection>
<intersection>10 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-39.5,-67.5,-39.5,-53.5</points>
<intersection>-67.5 9</intersection>
<intersection>-53.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-41,-67.5,-39.5,-67.5</points>
<connection>
<GID>130</GID>
<name>OUT_3</name></connection>
<intersection>-39.5 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>10,-48.5,11.5,-48.5</points>
<connection>
<GID>147</GID>
<name>IN_1</name></connection>
<intersection>10 0</intersection></hsegment></shape></wire>
<wire>
<ID>72 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-5.5,-59.5,-3.5,-59.5</points>
<connection>
<GID>145</GID>
<name>IN_1</name></connection>
<intersection>-5.5 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-5.5,-64.5,-5.5,-59.5</points>
<intersection>-64.5 15</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-38.5,-64.5,-3.5,-64.5</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>-38.5 17</intersection>
<intersection>-5.5 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>-38.5,-69.5,-38.5,-64.5</points>
<intersection>-69.5 18</intersection>
<intersection>-64.5 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>-41,-69.5,-38.5,-69.5</points>
<connection>
<GID>130</GID>
<name>OUT_2</name></connection>
<intersection>-38.5 17</intersection></hsegment></shape></wire>
<wire>
<ID>63 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4,-78.5,-4,-74.5</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<connection>
<GID>121</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>64 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-12,-84.5,-10,-84.5</points>
<connection>
<GID>137</GID>
<name>OUT</name></connection>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>-11.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-11.5,-84.5,-11.5,-79.5</points>
<intersection>-84.5 1</intersection>
<intersection>-79.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-11.5,-79.5,-10,-79.5</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>-11.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>3 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,-83,97.5,-83</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<connection>
<GID>15</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>78.5,-84,84,-84</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>78.5 4</intersection>
<intersection>81.5 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-84,78.5,-73</points>
<intersection>-84 2</intersection>
<intersection>-73 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>81.5,-89,81.5,-84</points>
<intersection>-89 15</intersection>
<intersection>-84 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>74.5,-73,78.5,-73</points>
<connection>
<GID>13</GID>
<name>OUT_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>81.5,-89,84,-89</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>81.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>1 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79.5,-82,84,-82</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>79.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>79.5,-87,79.5,-60</points>
<intersection>-87 16</intersection>
<intersection>-82 1</intersection>
<intersection>-60 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>74.5,-60,79.5,-60</points>
<connection>
<GID>8</GID>
<name>OUT_0</name></connection>
<intersection>79.5 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>79.5,-87,84,-87</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<intersection>79.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>57 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,-95.5,-24,-95.5</points>
<connection>
<GID>136</GID>
<name>IN_1</name></connection>
<intersection>-41 15</intersection>
<intersection>-30 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-30,-95.5,-30,-90.5</points>
<intersection>-95.5 1</intersection>
<intersection>-90.5 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-30,-90.5,-24,-90.5</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>-30 12</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>-41,-95.5,-41,-86.5</points>
<connection>
<GID>133</GID>
<name>OUT_0</name></connection>
<intersection>-95.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>77 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-40,-46.5,11.5,-46.5</points>
<connection>
<GID>147</GID>
<name>IN_0</name></connection>
<intersection>-40 6</intersection>
<intersection>9 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>9,-51.5,9,-46.5</points>
<intersection>-51.5 4</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>9,-51.5,11.5,-51.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>9 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-40,-54.5,-40,-46.5</points>
<intersection>-54.5 7</intersection>
<intersection>-46.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-41,-54.5,-40,-54.5</points>
<connection>
<GID>131</GID>
<name>OUT_3</name></connection>
<intersection>-40 6</intersection></hsegment></shape></wire>
<wire>
<ID>71 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-39,-57.5,-3.5,-57.5</points>
<connection>
<GID>145</GID>
<name>IN_0</name></connection>
<intersection>-39 18</intersection>
<intersection>-7.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-7.5,-62.5,-7.5,-57.5</points>
<intersection>-62.5 16</intersection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>-7.5,-62.5,-3.5,-62.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>-7.5 12</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>-39,-57.5,-39,-56.5</points>
<intersection>-57.5 1</intersection>
<intersection>-56.5 19</intersection></vsegment>
<hsegment>
<ID>19</ID>
<points>-41,-56.5,-39,-56.5</points>
<connection>
<GID>131</GID>
<name>OUT_2</name></connection>
<intersection>-39 18</intersection></hsegment></shape></wire>
<wire>
<ID>12 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-28.5,-6,-23,-6</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<connection>
<GID>70</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>55 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-25.5,-83.5,-18,-83.5</points>
<connection>
<GID>137</GID>
<name>IN_0</name></connection>
<connection>
<GID>129</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>54 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-37,-84.5,-31.5,-84.5</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>-37 4</intersection>
<intersection>-34 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-37,-84.5,-37,-73.5</points>
<intersection>-84.5 2</intersection>
<intersection>-73.5 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-34,-89.5,-34,-84.5</points>
<intersection>-89.5 15</intersection>
<intersection>-84.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>-41,-73.5,-37,-73.5</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>-37 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>-34,-89.5,-31.5,-89.5</points>
<connection>
<GID>128</GID>
<name>IN_1</name></connection>
<intersection>-34 11</intersection></hsegment></shape></wire>
<wire>
<ID>53 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-36,-82.5,-31.5,-82.5</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>-36 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>-36,-87.5,-36,-60.5</points>
<intersection>-87.5 16</intersection>
<intersection>-82.5 1</intersection>
<intersection>-60.5 15</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>-41,-60.5,-36,-60.5</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<intersection>-36 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>-36,-87.5,-31.5,-87.5</points>
<connection>
<GID>128</GID>
<name>IN_0</name></connection>
<intersection>-36 7</intersection></hsegment></shape></wire>
<wire>
<ID>11 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-25.5,-5,-25.5,1</points>
<intersection>-5 1</intersection>
<intersection>1 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-25.5,-5,-23,-5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>-25.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-28.5,1,-25.5,1</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>-25.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>5 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-41,2,-34.5,2</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>-39 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-39,-5,-39,2</points>
<intersection>-5 4</intersection>
<intersection>2 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-39,-5,-34.5,-5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>-39 3</intersection></hsegment></shape></wire>
<wire>
<ID>65 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-82.5,-11.5,-77.5</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>-82.5 23</intersection>
<intersection>-77.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-11.5,-77.5,-10,-77.5</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>-11.5,-82.5,-10,-82.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>-11.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>61 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-78.5,-19.5,-73.5</points>
<intersection>-78.5 2</intersection>
<intersection>-73.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-38,-78.5,-17.5,-78.5</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>-38 8</intersection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-19.5,-73.5,-17.5,-73.5</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>-38,-78.5,-38,-71.5</points>
<intersection>-78.5 2</intersection>
<intersection>-71.5 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>-41,-71.5,-38,-71.5</points>
<connection>
<GID>130</GID>
<name>OUT_1</name></connection>
<intersection>-38 8</intersection></hsegment></shape></wire>
<wire>
<ID>60 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20.5,-71.5,-17.5,-71.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>-20.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-20.5,-76.5,-20.5,-58.5</points>
<intersection>-76.5 4</intersection>
<intersection>-71.5 1</intersection>
<intersection>-58.5 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-20.5,-76.5,-17.5,-76.5</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>-20.5 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-41,-58.5,-20.5,-58.5</points>
<connection>
<GID>131</GID>
<name>OUT_1</name></connection>
<intersection>-20.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>6 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-37,-11,-37,0</points>
<intersection>-11 2</intersection>
<intersection>-7 3</intersection>
<intersection>0 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-37,0,-34.5,0</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>-37 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-41,-11,-37,-11</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>-37 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-37,-7,-34.5,-7</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>-37 0</intersection></hsegment></shape></wire>
<wire>
<ID>24 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>39.5,-8,39.5,0</points>
<intersection>-8 1</intersection>
<intersection>0 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>39.5,-8,42.5,-8</points>
<connection>
<GID>90</GID>
<name>IN_1</name></connection>
<intersection>39.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,0,39.5,0</points>
<connection>
<GID>89</GID>
<name>OUT</name></connection>
<intersection>39.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-7,30,-1</points>
<intersection>-7 2</intersection>
<intersection>-1 4</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>28.5,-7,30,-7</points>
<connection>
<GID>86</GID>
<name>OUT</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>30,-1,32,-1</points>
<connection>
<GID>89</GID>
<name>IN_1</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>19 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>18.5,1,32,1</points>
<connection>
<GID>79</GID>
<name>OUT</name></connection>
<connection>
<GID>89</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>84 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26,-73,26,-58.5</points>
<intersection>-73 1</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26,-73,36,-73</points>
<connection>
<GID>120</GID>
<name>IN_3</name></connection>
<intersection>26 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>25,-58.5,26,-58.5</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<intersection>26 0</intersection></hsegment></shape></wire>
<wire>
<ID>81 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>16,-59.5,19,-59.5</points>
<connection>
<GID>143</GID>
<name>OUT</name></connection>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>16.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>16.5,-59.5,16.5,-54.5</points>
<intersection>-59.5 1</intersection>
<intersection>-54.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>16.5,-54.5,19,-54.5</points>
<connection>
<GID>141</GID>
<name>IN_1</name></connection>
<intersection>16.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>82 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>17.5,-57.5,17.5,-52.5</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<intersection>-57.5 23</intersection>
<intersection>-52.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>17.5,-52.5,19,-52.5</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>17.5,-57.5,19,-57.5</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>17.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,-84,105.5,-84</points>
<connection>
<GID>21</GID>
<name>IN_1</name></connection>
<intersection>103.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>103.5,-84,103.5,-79</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>-84 1</intersection>
<intersection>-79 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>103.5,-79,105.5,-79</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>103.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>18 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-82,104,-77</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>-82 23</intersection>
<intersection>-77 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>104,-77,105.5,-77</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>104,-82,105.5,-82</points>
<connection>
<GID>21</GID>
<name>IN_0</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>27 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>89.5,-2.5,97,-2.5</points>
<connection>
<GID>100</GID>
<name>OUT</name></connection>
<connection>
<GID>92</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>30 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>89.5,-12.5,89.5,-7.5</points>
<intersection>-12.5 23</intersection>
<intersection>-7.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>89.5,-7.5,91,-7.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>89.5,-12.5,91,-12.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<intersection>89.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>78.5,-3.5,83.5,-3.5</points>
<connection>
<GID>100</GID>
<name>IN_1</name></connection>
<intersection>78.5 4</intersection>
<intersection>81.5 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-11,78.5,-3.5</points>
<intersection>-11 14</intersection>
<intersection>-3.5 2</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>81.5,-8.5,81.5,-3.5</points>
<intersection>-8.5 15</intersection>
<intersection>-3.5 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>74.5,-11,78.5,-11</points>
<connection>
<GID>99</GID>
<name>OUT_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>81.5,-8.5,83.5,-8.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>81.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>25 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>76.5,-1.5,83.5,-1.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>76.5 7</intersection>
<intersection>79.5 12</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>76.5,-1.5,76.5,2</points>
<intersection>-1.5 1</intersection>
<intersection>2 15</intersection></vsegment>
<vsegment>
<ID>12</ID>
<points>79.5,-6.5,79.5,-1.5</points>
<intersection>-6.5 16</intersection>
<intersection>-1.5 1</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>74.5,2,76.5,2</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<intersection>76.5 7</intersection></hsegment>
<hsegment>
<ID>16</ID>
<points>79.5,-6.5,83.5,-6.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>79.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>47 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,8.5,111,8.5</points>
<connection>
<GID>115</GID>
<name>OUT</name></connection>
<connection>
<GID>118</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>46 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,2.5,96,7.5</points>
<intersection>2.5 2</intersection>
<intersection>7.5 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>77.5,2.5,97.5,2.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>77.5 8</intersection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>96,7.5,97.5,7.5</points>
<connection>
<GID>115</GID>
<name>IN_1</name></connection>
<intersection>96 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>77.5,-9,77.5,2.5</points>
<intersection>-9 9</intersection>
<intersection>2.5 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>74.5,-9,77.5,-9</points>
<connection>
<GID>99</GID>
<name>OUT_1</name></connection>
<intersection>77.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>45 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95,9.5,97.5,9.5</points>
<connection>
<GID>115</GID>
<name>IN_0</name></connection>
<intersection>95 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>95,4,95,9.5</points>
<intersection>4 5</intersection>
<intersection>4.5 4</intersection>
<intersection>9.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>95,4.5,97.5,4.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>95 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>74.5,4,95,4</points>
<connection>
<GID>98</GID>
<name>OUT_1</name></connection>
<intersection>95 3</intersection></hsegment></shape></wire>
<wire>
<ID>48 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,2.5,111,6.5</points>
<connection>
<GID>116</GID>
<name>OUT</name></connection>
<connection>
<GID>118</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>51 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>115,-12.5,115,-2.5</points>
<intersection>-12.5 1</intersection>
<intersection>-2.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>115,-12.5,119,-12.5</points>
<connection>
<GID>91</GID>
<name>IN_1</name></connection>
<intersection>115 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111,-2.5,115,-2.5</points>
<connection>
<GID>117</GID>
<name>OUT</name></connection>
<intersection>115 0</intersection></hsegment></shape></wire>
<wire>
<ID>49 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103,-3.5,105,-3.5</points>
<connection>
<GID>117</GID>
<name>IN_1</name></connection>
<connection>
<GID>92</GID>
<name>OUT</name></connection>
<intersection>104 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>104,-3.5,104,1.5</points>
<intersection>-3.5 1</intersection>
<intersection>1.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>104,1.5,105,1.5</points>
<connection>
<GID>116</GID>
<name>IN_1</name></connection>
<intersection>104 3</intersection></hsegment></shape></wire>
<wire>
<ID>50 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>103.5,-1.5,103.5,3.5</points>
<connection>
<GID>114</GID>
<name>OUT</name></connection>
<intersection>-1.5 23</intersection>
<intersection>3.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>103.5,3.5,105,3.5</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<intersection>103.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>103.5,-1.5,105,-1.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>103.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-53,125.5,-48</points>
<intersection>-53 2</intersection>
<intersection>-48 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>76,-53,127,-53</points>
<connection>
<GID>23</GID>
<name>IN_1</name></connection>
<intersection>76 8</intersection>
<intersection>125.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>76,-67,76,-53</points>
<intersection>-67 9</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>74.5,-67,76,-67</points>
<connection>
<GID>13</GID>
<name>OUT_3</name></connection>
<intersection>76 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>125.5,-48,127,-48</points>
<connection>
<GID>22</GID>
<name>IN_1</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-46,127,-46</points>
<connection>
<GID>22</GID>
<name>IN_0</name></connection>
<intersection>75.5 6</intersection>
<intersection>124.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>124.5,-51,124.5,-46</points>
<intersection>-51 4</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>124.5,-51,127,-51</points>
<connection>
<GID>23</GID>
<name>IN_0</name></connection>
<intersection>124.5 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>75.5,-54,75.5,-46</points>
<intersection>-54 8</intersection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>74.5,-54,75.5,-54</points>
<connection>
<GID>8</GID>
<name>OUT_3</name></connection>
<intersection>75.5 6</intersection></hsegment></shape></wire>
<wire>
<ID>37 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-64,125.5,-60</points>
<connection>
<GID>25</GID>
<name>OUT</name></connection>
<connection>
<GID>26</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>36 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118,-58,125.5,-58</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<connection>
<GID>24</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>15 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-72,111.5,-72</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<connection>
<GID>19</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-78,96,-73</points>
<intersection>-78 2</intersection>
<intersection>-73 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-78,98,-78</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<intersection>77.5 8</intersection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>96,-73,98,-73</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>96 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>77.5,-78,77.5,-71</points>
<intersection>-78 2</intersection>
<intersection>-71 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>74.5,-71,77.5,-71</points>
<connection>
<GID>13</GID>
<name>OUT_1</name></connection>
<intersection>77.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>9 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95,-71,98,-71</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>95 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>95,-76,95,-58</points>
<intersection>-76 4</intersection>
<intersection>-71 1</intersection>
<intersection>-58 5</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>95,-76,98,-76</points>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>95 3</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>74.5,-58,95,-58</points>
<connection>
<GID>8</GID>
<name>OUT_1</name></connection>
<intersection>95 3</intersection></hsegment></shape></wire>
<wire>
<ID>42 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-47,140.5,-47</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<connection>
<GID>22</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>43 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,-53,140.5,-49</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<connection>
<GID>29</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>44 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131.5,-59,134.5,-59</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>131.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>131.5,-59,131.5,-54</points>
<intersection>-59 1</intersection>
<intersection>-54 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>131.5,-54,134.5,-54</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>131.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>59 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-57,133,-52</points>
<connection>
<GID>23</GID>
<name>OUT</name></connection>
<intersection>-57 23</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>133,-52,134.5,-52</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>133,-57,134.5,-57</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>38 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117.5,-70,119.5,-70</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>117.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>117.5,-73,117.5,-65</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>-70 1</intersection>
<intersection>-65 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>117.5,-65,119.5,-65</points>
<connection>
<GID>25</GID>
<name>IN_1</name></connection>
<intersection>117.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>39 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118,-68,118,-63</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>-68 23</intersection>
<intersection>-63 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>118,-63,119.5,-63</points>
<connection>
<GID>25</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>118,-68,119.5,-68</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>118 0</intersection></hsegment></shape></wire>
<wire>
<ID>35 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>110,-59,112,-59</points>
<connection>
<GID>24</GID>
<name>IN_1</name></connection>
<intersection>110 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>110,-64,110,-59</points>
<intersection>-64 15</intersection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>77,-64,112,-64</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>77 17</intersection>
<intersection>110 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>77,-69,77,-64</points>
<intersection>-69 18</intersection>
<intersection>-64 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>74.5,-69,77,-69</points>
<connection>
<GID>13</GID>
<name>OUT_2</name></connection>
<intersection>77 17</intersection></hsegment></shape></wire>
<wire>
<ID>34 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-56,112,-56</points>
<connection>
<GID>8</GID>
<name>OUT_2</name></connection>
<intersection>108 12</intersection>
<intersection>112 20</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>108,-62,108,-56</points>
<intersection>-62 16</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>108,-62,112,-62</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>108 12</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>112,-57,112,-56</points>
<connection>
<GID>24</GID>
<name>IN_0</name></connection>
<intersection>-56 1</intersection></vsegment></shape></wire>
<wire>
<ID>7 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-96.5,148,-96.5</points>
<intersection>88 12</intersection>
<intersection>91.5 19</intersection>
<intersection>148 15</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>88,-96.5,88,-90</points>
<intersection>-96.5 1</intersection>
<intersection>-90 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>88,-90,91.5,-90</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>88 12</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>148,-100,148,-96.5</points>
<intersection>-100 32</intersection>
<intersection>-96.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>91.5,-96.5,91.5,-95</points>
<connection>
<GID>14</GID>
<name>IN_1</name></connection>
<intersection>-96.5 1</intersection></vsegment>
<hsegment>
<ID>32</ID>
<points>146.5,-100,148,-100</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<intersection>148 15</intersection></hsegment></shape></wire>
<wire>
<ID>109 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>140.5,-105,140.5,-101</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<connection>
<GID>35</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>103 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-116,125.5,-112</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<connection>
<GID>38</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>105 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>118.5,-120,118.5,-115</points>
<intersection>-120 23</intersection>
<intersection>-115 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>118,-115,119.5,-115</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>118.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>118.5,-120,119.5,-120</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>118.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>102 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>118,-110,125.5,-110</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>108 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>133,-99,140.5,-99</points>
<connection>
<GID>41</GID>
<name>OUT</name></connection>
<connection>
<GID>35</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>110 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131.5,-111,134.5,-111</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>131.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>131.5,-111,131.5,-106</points>
<intersection>-111 1</intersection>
<intersection>-106 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>131.5,-106,134.5,-106</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<intersection>131.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>111 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-109,133,-104</points>
<connection>
<GID>40</GID>
<name>OUT</name></connection>
<intersection>-109 23</intersection>
<intersection>-104 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>133,-104,134.5,-104</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>133,-109,134.5,-109</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>133 0</intersection></hsegment></shape></wire>
<wire>
<ID>122 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-92,151,-58</points>
<intersection>-92 1</intersection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-92,174.5,-92</points>
<connection>
<GID>50</GID>
<name>IN_7</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140.5,-58,151,-58</points>
<connection>
<GID>4</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>121 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-93,150,-69</points>
<intersection>-93 1</intersection>
<intersection>-69 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,-93,174.5,-93</points>
<connection>
<GID>50</GID>
<name>IN_6</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125.5,-69,150,-69</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>120 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-94,149,-83</points>
<intersection>-94 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149,-94,174.5,-94</points>
<connection>
<GID>50</GID>
<name>IN_5</name></connection>
<intersection>149 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-83,149,-83</points>
<connection>
<GID>21</GID>
<name>OUT</name></connection>
<intersection>149 0</intersection></hsegment></shape></wire>
<wire>
<ID>119 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97.5,-95,174.5,-95</points>
<connection>
<GID>50</GID>
<name>IN_4</name></connection>
<intersection>97.5 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>97.5,-95,97.5,-94</points>
<connection>
<GID>14</GID>
<name>OUT</name></connection>
<intersection>-95 1</intersection></vsegment></shape></wire>
<wire>
<ID>118 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>149,-110,149,-96</points>
<intersection>-110 2</intersection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>149,-96,174.5,-96</points>
<connection>
<GID>50</GID>
<name>IN_3</name></connection>
<intersection>149 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>140.5,-110,149,-110</points>
<connection>
<GID>44</GID>
<name>OUT</name></connection>
<intersection>149 0</intersection></hsegment></shape></wire>
<wire>
<ID>117 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>150,-121,150,-97</points>
<intersection>-121 2</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>150,-97,174.5,-97</points>
<connection>
<GID>50</GID>
<name>IN_2</name></connection>
<intersection>150 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>125.5,-121,150,-121</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<intersection>150 0</intersection></hsegment></shape></wire>
<wire>
<ID>116 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>151,-135,151,-98</points>
<intersection>-135 2</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>151,-98,174.5,-98</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>151 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111.5,-135,151,-135</points>
<connection>
<GID>43</GID>
<name>OUT</name></connection>
<intersection>151 0</intersection></hsegment></shape></wire>
<wire>
<ID>104 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>117.5,-122,119.5,-122</points>
<connection>
<GID>33</GID>
<name>IN_1</name></connection>
<intersection>117.5 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>117.5,-125,117.5,-117</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>-122 1</intersection>
<intersection>-117 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>117.5,-117,119.5,-117</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>117.5 12</intersection></hsegment></shape></wire>
<wire>
<ID>94 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>104,-124,111.5,-124</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<connection>
<GID>36</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>89 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>97.5,-141,97.5,-137</points>
<connection>
<GID>53</GID>
<name>OUT</name></connection>
<connection>
<GID>55</GID>
<name>IN_1</name></connection></vsegment></shape></wire>
<wire>
<ID>88 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90,-135,97.5,-135</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<connection>
<GID>47</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>115 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,-146,152,-99</points>
<intersection>-146 2</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152,-99,174.5,-99</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>97.5,-146,152,-146</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire>
<wire>
<ID>90 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-147,91.5,-147</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>74.5 15</intersection>
<intersection>88 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>88,-147,88,-142</points>
<intersection>-147 1</intersection>
<intersection>-142 14</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>88,-142,91.5,-142</points>
<connection>
<GID>53</GID>
<name>IN_1</name></connection>
<intersection>88 12</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>74.5,-147,74.5,-138</points>
<connection>
<GID>48</GID>
<name>OUT_0</name></connection>
<intersection>-147 1</intersection></vsegment></shape></wire>
<wire>
<ID>91 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90,-145,90,-140</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>-145 23</intersection>
<intersection>-140 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>90,-140,91.5,-140</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>90,-145,91.5,-145</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>90 0</intersection></hsegment></shape></wire>
<wire>
<ID>95 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111.5,-130,111.5,-126</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<connection>
<GID>57</GID>
<name>OUT</name></connection></vsegment></shape></wire>
<wire>
<ID>96 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>103.5,-136,105.5,-136</points>
<connection>
<GID>55</GID>
<name>OUT</name></connection>
<connection>
<GID>43</GID>
<name>IN_1</name></connection>
<intersection>103.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>103.5,-136,103.5,-131</points>
<intersection>-136 1</intersection>
<intersection>-131 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>103.5,-131,105.5,-131</points>
<connection>
<GID>57</GID>
<name>IN_1</name></connection>
<intersection>103.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>97 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104.5,-134,104.5,-129</points>
<intersection>-134 23</intersection>
<intersection>-129 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>104,-129,105.5,-129</points>
<connection>
<GID>45</GID>
<name>OUT</name></connection>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment>
<hsegment>
<ID>23</ID>
<points>104.5,-134,105.5,-134</points>
<connection>
<GID>43</GID>
<name>IN_0</name></connection>
<intersection>104.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>125.5,-105,125.5,-100</points>
<intersection>-105 2</intersection>
<intersection>-100 10</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>76,-105,127,-105</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>76 8</intersection>
<intersection>125.5 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>76,-119,76,-105</points>
<intersection>-119 9</intersection>
<intersection>-105 2</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>74.5,-119,76,-119</points>
<connection>
<GID>58</GID>
<name>OUT_3</name></connection>
<intersection>76 8</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>125.5,-100,127,-100</points>
<connection>
<GID>41</GID>
<name>IN_1</name></connection>
<intersection>125.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>101 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>110,-111,112,-111</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<intersection>110 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>110,-116,110,-111</points>
<intersection>-116 15</intersection>
<intersection>-111 2</intersection></vsegment>
<hsegment>
<ID>15</ID>
<points>77,-116,112,-116</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<intersection>77 17</intersection>
<intersection>110 11</intersection></hsegment>
<vsegment>
<ID>17</ID>
<points>77,-121,77,-116</points>
<intersection>-121 18</intersection>
<intersection>-116 15</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>74.5,-121,77,-121</points>
<connection>
<GID>58</GID>
<name>OUT_2</name></connection>
<intersection>77 17</intersection></hsegment></shape></wire>
<wire>
<ID>93 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96,-130,96,-125</points>
<intersection>-130 2</intersection>
<intersection>-125 6</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>77.5,-130,98,-130</points>
<connection>
<GID>45</GID>
<name>IN_1</name></connection>
<intersection>77.5 8</intersection>
<intersection>96 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>96,-125,98,-125</points>
<connection>
<GID>36</GID>
<name>IN_1</name></connection>
<intersection>96 0</intersection></hsegment>
<vsegment>
<ID>8</ID>
<points>77.5,-130,77.5,-123</points>
<intersection>-130 2</intersection>
<intersection>-123 9</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>74.5,-123,77.5,-123</points>
<connection>
<GID>58</GID>
<name>OUT_1</name></connection>
<intersection>77.5 8</intersection></hsegment></shape></wire>
<wire>
<ID>87 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>78.5,-136,84,-136</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>78.5 4</intersection>
<intersection>81.5 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>78.5,-136,78.5,-125</points>
<intersection>-136 2</intersection>
<intersection>-125 14</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>81.5,-141,81.5,-136</points>
<intersection>-141 15</intersection>
<intersection>-136 2</intersection></vsegment>
<hsegment>
<ID>14</ID>
<points>74.5,-125,78.5,-125</points>
<connection>
<GID>58</GID>
<name>OUT_0</name></connection>
<intersection>78.5 4</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>81.5,-141,84,-141</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>81.5 11</intersection></hsegment></shape></wire>
<wire>
<ID>106 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>124,-98,127,-98</points>
<connection>
<GID>41</GID>
<name>IN_0</name></connection>
<intersection>124 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>124,-106,124,-98</points>
<intersection>-106 8</intersection>
<intersection>-103 4</intersection>
<intersection>-98 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>124,-103,127,-103</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>124 3</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>74.5,-106,124,-106</points>
<connection>
<GID>49</GID>
<name>OUT_3</name></connection>
<intersection>124 3</intersection></hsegment></shape></wire>
<wire>
<ID>100 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>77,-109,112,-109</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>77 20</intersection>
<intersection>108 12</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>108,-114,108,-109</points>
<intersection>-114 16</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>108,-114,112,-114</points>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>108 12</intersection></hsegment>
<vsegment>
<ID>20</ID>
<points>77,-109,77,-108</points>
<intersection>-109 1</intersection>
<intersection>-108 27</intersection></vsegment>
<hsegment>
<ID>27</ID>
<points>74.5,-108,77,-108</points>
<connection>
<GID>49</GID>
<name>OUT_2</name></connection>
<intersection>77 20</intersection></hsegment></shape></wire>
<wire>
<ID>92 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>78,-123,98,-123</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>78 6</intersection>
<intersection>95 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>95,-128,95,-123</points>
<intersection>-128 4</intersection>
<intersection>-123 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>95,-128,98,-128</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>95 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>78,-123,78,-110</points>
<intersection>-123 1</intersection>
<intersection>-110 13</intersection></vsegment>
<hsegment>
<ID>13</ID>
<points>74.5,-110,78,-110</points>
<connection>
<GID>49</GID>
<name>OUT_1</name></connection>
<intersection>78 6</intersection></hsegment></shape></wire>
<wire>
<ID>86 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79.5,-134,84,-134</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>79.5 7</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>79.5,-139,79.5,-112</points>
<intersection>-139 16</intersection>
<intersection>-134 1</intersection>
<intersection>-112 24</intersection></vsegment>
<hsegment>
<ID>16</ID>
<points>79.5,-139,84,-139</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>79.5 7</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>74.5,-112,79.5,-112</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>79.5 7</intersection></hsegment></shape></wire>
<wire>
<ID>123 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>152,-89.5,152,-48</points>
<intersection>-89.5 1</intersection>
<intersection>-48 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>152,-89.5,174.5,-89.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>152 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>146.5,-48,152,-48</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>152 0</intersection></hsegment></shape></wire></page 0></circuit>